module TX_FUNC__DOT__WR_PKT_PAYLOAD_10G(
MODE_10G,
MODE_1G,
MODE_2P5G,
MODE_5G,
RESETN,
TX_DATA,
TX_WE,
__START__,
clk,
rst,
__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__,
__ILA_TX_FUNC_valid__,
TXFIFO_BUFF_0,
TXFIFO_BUFF_1,
TXFIFO_BUFF_2,
TXFIFO_BUFF_3,
TXFIFO_BUFF_4,
TXFIFO_BUFF_5,
TXFIFO_BUFF_6,
TXFIFO_BUFF_7,
TXFIFO_BUFF_8,
TXFIFO_BUFF_9,
TXFIFO_BUFF_10,
TXFIFO_BUFF_11,
TXFIFO_BUFF_12,
TXFIFO_BUFF_13,
TXFIFO_BUFF_14,
TXFIFO_BUFF_15,
TXFIFO_BUFF_16,
TXFIFO_BUFF_17,
TXFIFO_BUFF_18,
TXFIFO_BUFF_19,
TXFIFO_BUFF_20,
TXFIFO_BUFF_21,
TXFIFO_BUFF_22,
TXFIFO_BUFF_23,
TXFIFO_BUFF_24,
TXFIFO_BUFF_25,
TXFIFO_BUFF_26,
TXFIFO_BUFF_27,
TXFIFO_BUFF_28,
TXFIFO_BUFF_29,
TXFIFO_BUFF_30,
TXFIFO_BUFF_31,
TXFIFO_FULL,
TXFIFO_WUSED_QWD,
TXFIFO_BUFF_RD_PTR,
TXFIFO_BUFF_WR_PTR,
TXFIFO_RD_OUTPUT,
TX_STATE,
TX_STATE_ENCAP,
TX_B2B_CNTR,
TX_PACKET_BYTE_CNT,
TX_WCNT,
XGMII_DOUT_REG,
XGMII_COUT_REG,
TX_PKT_SENT,
TX_BYTE_SENT,
CRC,
CRC_DAT_IN,
CRC_IN,
TX_WCNT_INI,
TX_BUF,
__COUNTER_start__n4
);
input            MODE_10G;
input            MODE_1G;
input            MODE_2P5G;
input            MODE_5G;
input            RESETN;
input     [63:0] TX_DATA;
input            TX_WE;
input            __START__;
input            clk;
input            rst;
output            __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__;
output            __ILA_TX_FUNC_valid__;
output     [63:0] TXFIFO_BUFF_0;
output     [63:0] TXFIFO_BUFF_1;
output     [63:0] TXFIFO_BUFF_2;
output     [63:0] TXFIFO_BUFF_3;
output     [63:0] TXFIFO_BUFF_4;
output     [63:0] TXFIFO_BUFF_5;
output     [63:0] TXFIFO_BUFF_6;
output     [63:0] TXFIFO_BUFF_7;
output     [63:0] TXFIFO_BUFF_8;
output     [63:0] TXFIFO_BUFF_9;
output     [63:0] TXFIFO_BUFF_10;
output     [63:0] TXFIFO_BUFF_11;
output     [63:0] TXFIFO_BUFF_12;
output     [63:0] TXFIFO_BUFF_13;
output     [63:0] TXFIFO_BUFF_14;
output     [63:0] TXFIFO_BUFF_15;
output     [63:0] TXFIFO_BUFF_16;
output     [63:0] TXFIFO_BUFF_17;
output     [63:0] TXFIFO_BUFF_18;
output     [63:0] TXFIFO_BUFF_19;
output     [63:0] TXFIFO_BUFF_20;
output     [63:0] TXFIFO_BUFF_21;
output     [63:0] TXFIFO_BUFF_22;
output     [63:0] TXFIFO_BUFF_23;
output     [63:0] TXFIFO_BUFF_24;
output     [63:0] TXFIFO_BUFF_25;
output     [63:0] TXFIFO_BUFF_26;
output     [63:0] TXFIFO_BUFF_27;
output     [63:0] TXFIFO_BUFF_28;
output     [63:0] TXFIFO_BUFF_29;
output     [63:0] TXFIFO_BUFF_30;
output     [63:0] TXFIFO_BUFF_31;
output reg            TXFIFO_FULL;
output reg     [12:0] TXFIFO_WUSED_QWD;
output reg      [4:0] TXFIFO_BUFF_RD_PTR;
output reg      [4:0] TXFIFO_BUFF_WR_PTR;
output reg     [63:0] TXFIFO_RD_OUTPUT;
output reg      [4:0] TX_STATE;
output reg      [7:0] TX_STATE_ENCAP;
output reg      [5:0] TX_B2B_CNTR;
output reg     [15:0] TX_PACKET_BYTE_CNT;
output reg     [15:0] TX_WCNT;
output reg     [63:0] XGMII_DOUT_REG;
output reg      [7:0] XGMII_COUT_REG;
output reg     [31:0] TX_PKT_SENT;
output reg     [31:0] TX_BYTE_SENT;
output reg     [31:0] CRC;
output reg     [63:0] CRC_DAT_IN;
output reg     [31:0] CRC_IN;
output reg     [15:0] TX_WCNT_INI;
output reg     [63:0] TX_BUF;
output reg      [7:0] __COUNTER_start__n4;
(* keep *) wire     [63:0] CRC_DAT_IN_randinit;
(* keep *) wire     [31:0] CRC_IN_randinit;
(* keep *) wire     [31:0] CRC_randinit;
wire            MODE_10G;
wire            MODE_1G;
wire            MODE_2P5G;
wire            MODE_5G;
wire            RESETN;
wire     [63:0] TXFIFO_BUFF_0;
wire     [63:0] TXFIFO_BUFF_1;
wire     [63:0] TXFIFO_BUFF_10;
wire     [63:0] TXFIFO_BUFF_11;
wire     [63:0] TXFIFO_BUFF_12;
wire     [63:0] TXFIFO_BUFF_13;
wire     [63:0] TXFIFO_BUFF_14;
wire     [63:0] TXFIFO_BUFF_15;
wire     [63:0] TXFIFO_BUFF_16;
wire     [63:0] TXFIFO_BUFF_17;
wire     [63:0] TXFIFO_BUFF_18;
wire     [63:0] TXFIFO_BUFF_19;
wire     [63:0] TXFIFO_BUFF_2;
wire     [63:0] TXFIFO_BUFF_20;
wire     [63:0] TXFIFO_BUFF_21;
wire     [63:0] TXFIFO_BUFF_22;
wire     [63:0] TXFIFO_BUFF_23;
wire     [63:0] TXFIFO_BUFF_24;
wire     [63:0] TXFIFO_BUFF_25;
wire     [63:0] TXFIFO_BUFF_26;
wire     [63:0] TXFIFO_BUFF_27;
wire     [63:0] TXFIFO_BUFF_28;
wire     [63:0] TXFIFO_BUFF_29;
wire     [63:0] TXFIFO_BUFF_3;
wire     [63:0] TXFIFO_BUFF_30;
wire     [63:0] TXFIFO_BUFF_31;
wire     [63:0] TXFIFO_BUFF_4;
wire     [63:0] TXFIFO_BUFF_5;
wire     [63:0] TXFIFO_BUFF_6;
wire     [63:0] TXFIFO_BUFF_7;
wire     [63:0] TXFIFO_BUFF_8;
wire     [63:0] TXFIFO_BUFF_9;
(* keep *) wire      [4:0] TXFIFO_BUFF_RD_PTR_randinit;
(* keep *) wire      [4:0] TXFIFO_BUFF_WR_PTR_randinit;
(* keep *) wire            TXFIFO_FULL_randinit;
(* keep *) wire     [63:0] TXFIFO_RD_OUTPUT_randinit;
(* keep *) wire     [12:0] TXFIFO_WUSED_QWD_randinit;
(* keep *) wire      [5:0] TX_B2B_CNTR_randinit;
(* keep *) wire     [63:0] TX_BUF_randinit;
(* keep *) wire     [31:0] TX_BYTE_SENT_randinit;
wire     [63:0] TX_DATA;
(* keep *) wire     [15:0] TX_PACKET_BYTE_CNT_randinit;
(* keep *) wire     [31:0] TX_PKT_SENT_randinit;
(* keep *) wire      [7:0] TX_STATE_ENCAP_randinit;
(* keep *) wire      [4:0] TX_STATE_randinit;
(* keep *) wire     [15:0] TX_WCNT_INI_randinit;
(* keep *) wire     [15:0] TX_WCNT_randinit;
wire            TX_WE;
(* keep *) wire      [7:0] XGMII_COUT_REG_randinit;
(* keep *) wire     [63:0] XGMII_DOUT_REG_randinit;
wire            __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__;
wire            __ILA_TX_FUNC_valid__;
wire            __START__;
wire            clk;
wire            n0____DOLLAR__124;
wire     [63:0] n100____DOLLAR__3086;
wire     [63:0] n101____DOLLAR__3091;
wire     [63:0] n102____DOLLAR__3096;
wire     [63:0] n103____DOLLAR__3101;
wire     [63:0] n104____DOLLAR__3065;
wire     [63:0] n105____DOLLAR__3106;
wire     [63:0] n106____DOLLAR__3149;
wire     [63:0] n107____DOLLAR__3154;
wire            n108____DOLLAR__2865;
wire            n109____DOLLAR__2855;
wire      [4:0] n10____DOLLAR__486;
wire            n110____DOLLAR__2857;
wire            n111____DOLLAR__2859;
wire            n112____DOLLAR__2850;
wire            n113____DOLLAR__2843;
wire            n114____DOLLAR__2836;
wire            n115____DOLLAR__2829;
wire            n116____DOLLAR__2822;
wire            n117____DOLLAR__2815;
wire            n118____DOLLAR__2808;
wire      [7:0] n119____DOLLAR__2810;
wire      [4:0] n11____DOLLAR__493;
wire      [7:0] n120____DOLLAR__2817;
wire      [7:0] n121____DOLLAR__2824;
wire      [7:0] n122____DOLLAR__2831;
wire      [7:0] n123____DOLLAR__2838;
wire      [7:0] n124____DOLLAR__2845;
wire      [7:0] n125____DOLLAR__2852;
wire            n126____DOLLAR__2799;
wire            n127____DOLLAR__2794;
wire            n128____DOLLAR__2787;
wire            n129____DOLLAR__2780;
wire      [4:0] n12____DOLLAR__498;
wire            n130____DOLLAR__2773;
wire            n131____DOLLAR__2766;
wire            n132____DOLLAR__2759;
wire            n133____DOLLAR__2752;
wire      [7:0] n134____DOLLAR__2754;
wire      [7:0] n135____DOLLAR__2761;
wire      [7:0] n136____DOLLAR__2768;
wire      [7:0] n137____DOLLAR__2775;
wire      [7:0] n138____DOLLAR__2782;
wire      [7:0] n139____DOLLAR__2789;
wire            n13____DOLLAR__481;
wire      [7:0] n140____DOLLAR__2796;
wire      [7:0] n141____DOLLAR__2801;
wire      [7:0] n142____DOLLAR__2860;
wire      [7:0] n143____DOLLAR__2867;
wire            n144____DOLLAR__2705;
wire     [31:0] n145____DOLLAR__2696;
wire     [31:0] n146____DOLLAR__2697;
wire     [31:0] n147____DOLLAR__2690;
wire     [31:0] n148____DOLLAR__2691;
wire     [31:0] n149____DOLLAR__2698;
wire     [63:0] n14____DOLLAR__477;
wire     [31:0] n150____DOLLAR__2684;
wire     [31:0] n151____DOLLAR__2685;
wire     [31:0] n152____DOLLAR__2699;
wire     [31:0] n153____DOLLAR__2678;
wire     [31:0] n154____DOLLAR__2674;
wire     [31:0] n155____DOLLAR__2679;
wire     [31:0] n156____DOLLAR__2700;
wire     [31:0] n157____DOLLAR__2701;
wire     [31:0] n158____DOLLAR__2707;
wire            n159____DOLLAR__508;
wire     [63:0] n15____DOLLAR__483;
wire            n160____DOLLAR__743;
wire            n161____DOLLAR__738;
wire      [7:0] n162____DOLLAR__728;
wire     [55:0] n163____DOLLAR__726;
wire     [63:0] n164____DOLLAR__734;
wire            n165____DOLLAR__715;
wire     [15:0] n166____DOLLAR__705;
wire     [47:0] n167____DOLLAR__703;
wire     [63:0] n168____DOLLAR__711;
wire            n169____DOLLAR__692;
wire            n16____DOLLAR__3169;
wire     [23:0] n170____DOLLAR__682;
wire     [39:0] n171____DOLLAR__680;
wire     [63:0] n172____DOLLAR__688;
wire            n173____DOLLAR__669;
wire     [31:0] n174____DOLLAR__659;
wire     [63:0] n175____DOLLAR__665;
wire            n176____DOLLAR__654;
wire     [39:0] n177____DOLLAR__644;
wire     [63:0] n178____DOLLAR__650;
wire            n179____DOLLAR__639;
wire      [4:0] n17____DOLLAR__3171;
wire     [47:0] n180____DOLLAR__629;
wire     [63:0] n181____DOLLAR__635;
wire     [55:0] n182____DOLLAR__619;
wire     [63:0] n183____DOLLAR__625;
wire     [63:0] n184____DOLLAR__641;
wire     [63:0] n185____DOLLAR__656;
wire     [63:0] n186____DOLLAR__671;
wire     [63:0] n187____DOLLAR__694;
wire     [63:0] n188____DOLLAR__717;
wire     [63:0] n189____DOLLAR__740;
wire            n18____DOLLAR__3176;
wire     [63:0] n190____DOLLAR__745;
wire            n191____DOLLAR__614;
wire            n192____DOLLAR__609;
wire      [7:0] n193____DOLLAR__599;
wire     [55:0] n194____DOLLAR__597;
wire     [63:0] n195____DOLLAR__605;
wire            n196____DOLLAR__594;
wire     [15:0] n197____DOLLAR__584;
wire     [47:0] n198____DOLLAR__582;
wire     [63:0] n199____DOLLAR__590;
wire      [7:0] n19____DOLLAR__3178;
wire            n1____DOLLAR__467;
wire            n200____DOLLAR__579;
wire     [23:0] n201____DOLLAR__569;
wire     [39:0] n202____DOLLAR__567;
wire     [63:0] n203____DOLLAR__575;
wire            n204____DOLLAR__564;
wire     [31:0] n205____DOLLAR__554;
wire     [31:0] n206____DOLLAR__552;
wire     [63:0] n207____DOLLAR__560;
wire            n208____DOLLAR__549;
wire     [39:0] n209____DOLLAR__539;
wire            n20____DOLLAR__3160;
wire     [23:0] n210____DOLLAR__537;
wire     [63:0] n211____DOLLAR__545;
wire            n212____DOLLAR__534;
wire     [47:0] n213____DOLLAR__524;
wire     [15:0] n214____DOLLAR__522;
wire     [63:0] n215____DOLLAR__530;
wire     [55:0] n216____DOLLAR__514;
wire      [7:0] n217____DOLLAR__512;
wire     [63:0] n218____DOLLAR__520;
wire     [63:0] n219____DOLLAR__536;
wire      [5:0] n21____DOLLAR__3157;
wire     [63:0] n220____DOLLAR__551;
wire     [63:0] n221____DOLLAR__566;
wire     [63:0] n222____DOLLAR__581;
wire     [63:0] n223____DOLLAR__596;
wire     [63:0] n224____DOLLAR__611;
wire     [63:0] n225____DOLLAR__616;
wire     [63:0] n226____DOLLAR__746;
wire            n227____DOLLAR__2663;
wire      [7:0] n228____DOLLAR__756;
wire      [7:0] n229____DOLLAR__749;
wire      [5:0] n22____DOLLAR__3162;
wire      [7:0] n230____DOLLAR__758;
wire      [7:0] n231____DOLLAR__759;
wire            n232____DOLLAR__864;
wire            n233____DOLLAR__857;
wire            n234____DOLLAR__850;
wire            n235____DOLLAR__843;
wire            n236____DOLLAR__836;
wire            n237____DOLLAR__829;
wire            n238____DOLLAR__822;
wire            n239____DOLLAR__815;
wire     [15:0] n23____DOLLAR__3181;
wire            n240____DOLLAR__808;
wire            n241____DOLLAR__801;
wire            n242____DOLLAR__794;
wire            n243____DOLLAR__787;
wire            n244____DOLLAR__780;
wire            n245____DOLLAR__773;
wire            n246____DOLLAR__766;
wire     [31:0] n247____DOLLAR__768;
wire     [31:0] n248____DOLLAR__775;
wire     [31:0] n249____DOLLAR__782;
wire            n24____DOLLAR__3152;
wire     [31:0] n250____DOLLAR__789;
wire     [31:0] n251____DOLLAR__796;
wire     [31:0] n252____DOLLAR__803;
wire     [31:0] n253____DOLLAR__810;
wire     [31:0] n254____DOLLAR__817;
wire     [31:0] n255____DOLLAR__824;
wire     [31:0] n256____DOLLAR__831;
wire     [31:0] n257____DOLLAR__838;
wire     [31:0] n258____DOLLAR__845;
wire     [31:0] n259____DOLLAR__852;
wire            n25____DOLLAR__3144;
wire     [31:0] n260____DOLLAR__859;
wire     [31:0] n261____DOLLAR__866;
wire     [31:0] n262____DOLLAR__753;
wire     [31:0] n263____DOLLAR__867;
wire      [7:0] n264____DOLLAR__876;
wire      [7:0] n265____DOLLAR__875;
wire      [7:0] n266____DOLLAR__878;
wire      [7:0] n267____DOLLAR__879;
wire            n268____DOLLAR__984;
wire            n269____DOLLAR__977;
wire            n26____DOLLAR__3146;
wire            n270____DOLLAR__970;
wire            n271____DOLLAR__963;
wire            n272____DOLLAR__956;
wire            n273____DOLLAR__949;
wire            n274____DOLLAR__942;
wire            n275____DOLLAR__935;
wire            n276____DOLLAR__928;
wire            n277____DOLLAR__921;
wire            n278____DOLLAR__914;
wire            n279____DOLLAR__907;
wire            n27____DOLLAR__3148;
wire            n280____DOLLAR__900;
wire            n281____DOLLAR__893;
wire            n282____DOLLAR__886;
wire     [31:0] n283____DOLLAR__888;
wire     [31:0] n284____DOLLAR__895;
wire     [31:0] n285____DOLLAR__902;
wire     [31:0] n286____DOLLAR__909;
wire     [31:0] n287____DOLLAR__916;
wire     [31:0] n288____DOLLAR__923;
wire     [31:0] n289____DOLLAR__930;
wire      [2:0] n28____DOLLAR__510;
wire     [31:0] n290____DOLLAR__937;
wire     [31:0] n291____DOLLAR__944;
wire     [31:0] n292____DOLLAR__951;
wire     [31:0] n293____DOLLAR__958;
wire     [31:0] n294____DOLLAR__965;
wire     [31:0] n295____DOLLAR__972;
wire     [31:0] n296____DOLLAR__979;
wire     [31:0] n297____DOLLAR__986;
wire     [31:0] n298____DOLLAR__870;
wire     [31:0] n299____DOLLAR__987;
wire            n29____DOLLAR__3139;
wire            n2____DOLLAR__472;
wire      [7:0] n300____DOLLAR__995;
wire      [7:0] n301____DOLLAR__988;
wire      [7:0] n302____DOLLAR__997;
wire      [7:0] n303____DOLLAR__998;
wire            n304____DOLLAR__1103;
wire            n305____DOLLAR__1096;
wire            n306____DOLLAR__1089;
wire            n307____DOLLAR__1082;
wire            n308____DOLLAR__1075;
wire            n309____DOLLAR__1068;
wire            n30____DOLLAR__3134;
wire            n310____DOLLAR__1061;
wire            n311____DOLLAR__1054;
wire            n312____DOLLAR__1047;
wire            n313____DOLLAR__1040;
wire            n314____DOLLAR__1033;
wire            n315____DOLLAR__1026;
wire            n316____DOLLAR__1019;
wire            n317____DOLLAR__1012;
wire            n318____DOLLAR__1005;
wire     [31:0] n319____DOLLAR__1007;
wire     [31:0] n31____DOLLAR__2739;
wire     [31:0] n320____DOLLAR__1014;
wire     [31:0] n321____DOLLAR__1021;
wire     [31:0] n322____DOLLAR__1028;
wire     [31:0] n323____DOLLAR__1035;
wire     [31:0] n324____DOLLAR__1042;
wire     [31:0] n325____DOLLAR__1049;
wire     [31:0] n326____DOLLAR__1056;
wire     [31:0] n327____DOLLAR__1063;
wire     [31:0] n328____DOLLAR__1070;
wire     [31:0] n329____DOLLAR__1077;
wire     [31:0] n32____DOLLAR__2740;
wire     [31:0] n330____DOLLAR__1084;
wire     [31:0] n331____DOLLAR__1091;
wire     [31:0] n332____DOLLAR__1098;
wire     [31:0] n333____DOLLAR__1105;
wire     [31:0] n334____DOLLAR__992;
wire     [31:0] n335____DOLLAR__1106;
wire      [7:0] n336____DOLLAR__1115;
wire      [7:0] n337____DOLLAR__1114;
wire      [7:0] n338____DOLLAR__1117;
wire      [7:0] n339____DOLLAR__1118;
wire     [31:0] n33____DOLLAR__2733;
wire            n340____DOLLAR__1223;
wire            n341____DOLLAR__1216;
wire            n342____DOLLAR__1209;
wire            n343____DOLLAR__1202;
wire            n344____DOLLAR__1195;
wire            n345____DOLLAR__1188;
wire            n346____DOLLAR__1181;
wire            n347____DOLLAR__1174;
wire            n348____DOLLAR__1167;
wire            n349____DOLLAR__1160;
wire     [31:0] n34____DOLLAR__2734;
wire            n350____DOLLAR__1153;
wire            n351____DOLLAR__1146;
wire            n352____DOLLAR__1139;
wire            n353____DOLLAR__1132;
wire            n354____DOLLAR__1125;
wire     [31:0] n355____DOLLAR__1127;
wire     [31:0] n356____DOLLAR__1134;
wire     [31:0] n357____DOLLAR__1141;
wire     [31:0] n358____DOLLAR__1148;
wire     [31:0] n359____DOLLAR__1155;
wire     [31:0] n35____DOLLAR__2741;
wire     [31:0] n360____DOLLAR__1162;
wire     [31:0] n361____DOLLAR__1169;
wire     [31:0] n362____DOLLAR__1176;
wire     [31:0] n363____DOLLAR__1183;
wire     [31:0] n364____DOLLAR__1190;
wire     [31:0] n365____DOLLAR__1197;
wire     [31:0] n366____DOLLAR__1204;
wire     [31:0] n367____DOLLAR__1211;
wire     [31:0] n368____DOLLAR__1218;
wire     [31:0] n369____DOLLAR__1225;
wire     [31:0] n36____DOLLAR__2727;
wire     [31:0] n370____DOLLAR__1109;
wire     [31:0] n371____DOLLAR__1226;
wire      [7:0] n372____DOLLAR__1234;
wire      [7:0] n373____DOLLAR__1227;
wire      [7:0] n374____DOLLAR__1236;
wire      [7:0] n375____DOLLAR__1237;
wire            n376____DOLLAR__1342;
wire            n377____DOLLAR__1335;
wire            n378____DOLLAR__1328;
wire            n379____DOLLAR__1321;
wire     [31:0] n37____DOLLAR__2728;
wire            n380____DOLLAR__1314;
wire            n381____DOLLAR__1307;
wire            n382____DOLLAR__1300;
wire            n383____DOLLAR__1293;
wire            n384____DOLLAR__1286;
wire            n385____DOLLAR__1279;
wire            n386____DOLLAR__1272;
wire            n387____DOLLAR__1265;
wire            n388____DOLLAR__1258;
wire            n389____DOLLAR__1251;
wire     [31:0] n38____DOLLAR__2742;
wire            n390____DOLLAR__1244;
wire     [31:0] n391____DOLLAR__1246;
wire     [31:0] n392____DOLLAR__1253;
wire     [31:0] n393____DOLLAR__1260;
wire     [31:0] n394____DOLLAR__1267;
wire     [31:0] n395____DOLLAR__1274;
wire     [31:0] n396____DOLLAR__1281;
wire     [31:0] n397____DOLLAR__1288;
wire     [31:0] n398____DOLLAR__1295;
wire     [31:0] n399____DOLLAR__1302;
wire     [31:0] n39____DOLLAR__2721;
wire            n3____DOLLAR__474;
wire     [31:0] n400____DOLLAR__1309;
wire     [31:0] n401____DOLLAR__1316;
wire     [31:0] n402____DOLLAR__1323;
wire     [31:0] n403____DOLLAR__1330;
wire     [31:0] n404____DOLLAR__1337;
wire     [31:0] n405____DOLLAR__1344;
wire     [31:0] n406____DOLLAR__1231;
wire     [31:0] n407____DOLLAR__1345;
wire      [7:0] n408____DOLLAR__1354;
wire      [7:0] n409____DOLLAR__1353;
wire     [31:0] n40____DOLLAR__2717;
wire      [7:0] n410____DOLLAR__1356;
wire      [7:0] n411____DOLLAR__1357;
wire            n412____DOLLAR__1462;
wire            n413____DOLLAR__1455;
wire            n414____DOLLAR__1448;
wire            n415____DOLLAR__1441;
wire            n416____DOLLAR__1434;
wire            n417____DOLLAR__1427;
wire            n418____DOLLAR__1420;
wire            n419____DOLLAR__1413;
wire     [31:0] n41____DOLLAR__2722;
wire            n420____DOLLAR__1406;
wire            n421____DOLLAR__1399;
wire            n422____DOLLAR__1392;
wire            n423____DOLLAR__1385;
wire            n424____DOLLAR__1378;
wire            n425____DOLLAR__1371;
wire            n426____DOLLAR__1364;
wire     [31:0] n427____DOLLAR__1366;
wire     [31:0] n428____DOLLAR__1373;
wire     [31:0] n429____DOLLAR__1380;
wire     [31:0] n42____DOLLAR__2743;
wire     [31:0] n430____DOLLAR__1387;
wire     [31:0] n431____DOLLAR__1394;
wire     [31:0] n432____DOLLAR__1401;
wire     [31:0] n433____DOLLAR__1408;
wire     [31:0] n434____DOLLAR__1415;
wire     [31:0] n435____DOLLAR__1422;
wire     [31:0] n436____DOLLAR__1429;
wire     [31:0] n437____DOLLAR__1436;
wire     [31:0] n438____DOLLAR__1443;
wire     [31:0] n439____DOLLAR__1450;
wire      [7:0] n43____DOLLAR__2869;
wire     [31:0] n440____DOLLAR__1457;
wire     [31:0] n441____DOLLAR__1464;
wire     [31:0] n442____DOLLAR__1348;
wire     [31:0] n443____DOLLAR__1465;
wire      [7:0] n444____DOLLAR__1473;
wire      [7:0] n445____DOLLAR__1466;
wire      [7:0] n446____DOLLAR__1475;
wire      [7:0] n447____DOLLAR__1476;
wire            n448____DOLLAR__1581;
wire            n449____DOLLAR__1574;
wire     [39:0] n44____DOLLAR__2875;
wire            n450____DOLLAR__1567;
wire            n451____DOLLAR__1560;
wire            n452____DOLLAR__1553;
wire            n453____DOLLAR__1546;
wire            n454____DOLLAR__1539;
wire            n455____DOLLAR__1532;
wire            n456____DOLLAR__1525;
wire            n457____DOLLAR__1518;
wire            n458____DOLLAR__1511;
wire            n459____DOLLAR__1504;
wire     [63:0] n45____DOLLAR__2883;
wire            n460____DOLLAR__1497;
wire            n461____DOLLAR__1490;
wire            n462____DOLLAR__1483;
wire     [31:0] n463____DOLLAR__1485;
wire     [31:0] n464____DOLLAR__1492;
wire     [31:0] n465____DOLLAR__1499;
wire     [31:0] n466____DOLLAR__1506;
wire     [31:0] n467____DOLLAR__1513;
wire     [31:0] n468____DOLLAR__1520;
wire     [31:0] n469____DOLLAR__1527;
wire            n46____DOLLAR__3129;
wire     [31:0] n470____DOLLAR__1534;
wire     [31:0] n471____DOLLAR__1541;
wire     [31:0] n472____DOLLAR__1548;
wire     [31:0] n473____DOLLAR__1555;
wire     [31:0] n474____DOLLAR__1562;
wire     [31:0] n475____DOLLAR__1569;
wire     [31:0] n476____DOLLAR__1576;
wire     [31:0] n477____DOLLAR__1583;
wire     [31:0] n478____DOLLAR__1470;
wire     [31:0] n479____DOLLAR__1584;
wire     [15:0] n47____DOLLAR__2885;
wire      [7:0] n480____DOLLAR__1593;
wire      [7:0] n481____DOLLAR__1592;
wire      [7:0] n482____DOLLAR__1595;
wire      [7:0] n483____DOLLAR__1596;
wire            n484____DOLLAR__1701;
wire            n485____DOLLAR__1694;
wire            n486____DOLLAR__1687;
wire            n487____DOLLAR__1680;
wire            n488____DOLLAR__1673;
wire            n489____DOLLAR__1666;
wire     [47:0] n48____DOLLAR__2891;
wire            n490____DOLLAR__1659;
wire            n491____DOLLAR__1652;
wire            n492____DOLLAR__1645;
wire            n493____DOLLAR__1638;
wire            n494____DOLLAR__1631;
wire            n495____DOLLAR__1624;
wire            n496____DOLLAR__1617;
wire            n497____DOLLAR__1610;
wire            n498____DOLLAR__1603;
wire     [31:0] n499____DOLLAR__1605;
wire     [63:0] n49____DOLLAR__2899;
wire     [31:0] n500____DOLLAR__1612;
wire     [31:0] n501____DOLLAR__1619;
wire     [31:0] n502____DOLLAR__1626;
wire     [31:0] n503____DOLLAR__1633;
wire     [31:0] n504____DOLLAR__1640;
wire     [31:0] n505____DOLLAR__1647;
wire     [31:0] n506____DOLLAR__1654;
wire     [31:0] n507____DOLLAR__1661;
wire     [31:0] n508____DOLLAR__1668;
wire     [31:0] n509____DOLLAR__1675;
wire            n50____DOLLAR__3124;
wire     [31:0] n510____DOLLAR__1682;
wire     [31:0] n511____DOLLAR__1689;
wire     [31:0] n512____DOLLAR__1696;
wire     [31:0] n513____DOLLAR__1703;
wire     [31:0] n514____DOLLAR__1587;
wire     [31:0] n515____DOLLAR__1704;
wire      [7:0] n516____DOLLAR__1712;
wire      [7:0] n517____DOLLAR__1705;
wire      [7:0] n518____DOLLAR__1714;
wire      [7:0] n519____DOLLAR__1715;
wire     [23:0] n51____DOLLAR__2901;
wire            n520____DOLLAR__1820;
wire            n521____DOLLAR__1813;
wire            n522____DOLLAR__1806;
wire            n523____DOLLAR__1799;
wire            n524____DOLLAR__1792;
wire            n525____DOLLAR__1785;
wire            n526____DOLLAR__1778;
wire            n527____DOLLAR__1771;
wire            n528____DOLLAR__1764;
wire            n529____DOLLAR__1757;
wire     [55:0] n52____DOLLAR__2907;
wire            n530____DOLLAR__1750;
wire            n531____DOLLAR__1743;
wire            n532____DOLLAR__1736;
wire            n533____DOLLAR__1729;
wire            n534____DOLLAR__1722;
wire     [31:0] n535____DOLLAR__1724;
wire     [31:0] n536____DOLLAR__1731;
wire     [31:0] n537____DOLLAR__1738;
wire     [31:0] n538____DOLLAR__1745;
wire     [31:0] n539____DOLLAR__1752;
wire     [63:0] n53____DOLLAR__2915;
wire     [31:0] n540____DOLLAR__1759;
wire     [31:0] n541____DOLLAR__1766;
wire     [31:0] n542____DOLLAR__1773;
wire     [31:0] n543____DOLLAR__1780;
wire     [31:0] n544____DOLLAR__1787;
wire     [31:0] n545____DOLLAR__1794;
wire     [31:0] n546____DOLLAR__1801;
wire     [31:0] n547____DOLLAR__1808;
wire     [31:0] n548____DOLLAR__1815;
wire     [31:0] n549____DOLLAR__1822;
wire            n54____DOLLAR__3119;
wire     [31:0] n550____DOLLAR__1709;
wire     [31:0] n551____DOLLAR__1823;
wire      [7:0] n552____DOLLAR__1832;
wire      [7:0] n553____DOLLAR__1831;
wire      [7:0] n554____DOLLAR__1834;
wire      [7:0] n555____DOLLAR__1835;
wire            n556____DOLLAR__1940;
wire            n557____DOLLAR__1933;
wire            n558____DOLLAR__1926;
wire            n559____DOLLAR__1919;
wire     [31:0] n55____DOLLAR__2917;
wire            n560____DOLLAR__1912;
wire            n561____DOLLAR__1905;
wire            n562____DOLLAR__1898;
wire            n563____DOLLAR__1891;
wire            n564____DOLLAR__1884;
wire            n565____DOLLAR__1877;
wire            n566____DOLLAR__1870;
wire            n567____DOLLAR__1863;
wire            n568____DOLLAR__1856;
wire            n569____DOLLAR__1849;
wire     [63:0] n56____DOLLAR__2923;
wire            n570____DOLLAR__1842;
wire     [31:0] n571____DOLLAR__1844;
wire     [31:0] n572____DOLLAR__1851;
wire     [31:0] n573____DOLLAR__1858;
wire     [31:0] n574____DOLLAR__1865;
wire     [31:0] n575____DOLLAR__1872;
wire     [31:0] n576____DOLLAR__1879;
wire     [31:0] n577____DOLLAR__1886;
wire     [31:0] n578____DOLLAR__1893;
wire     [31:0] n579____DOLLAR__1900;
wire            n57____DOLLAR__3114;
wire     [31:0] n580____DOLLAR__1907;
wire     [31:0] n581____DOLLAR__1914;
wire     [31:0] n582____DOLLAR__1921;
wire     [31:0] n583____DOLLAR__1928;
wire     [31:0] n584____DOLLAR__1935;
wire     [31:0] n585____DOLLAR__1942;
wire     [31:0] n586____DOLLAR__1826;
wire     [31:0] n587____DOLLAR__1943;
wire      [7:0] n588____DOLLAR__1951;
wire      [7:0] n589____DOLLAR__1944;
wire     [23:0] n58____DOLLAR__2927;
wire      [7:0] n590____DOLLAR__1953;
wire      [7:0] n591____DOLLAR__1954;
wire            n592____DOLLAR__2059;
wire            n593____DOLLAR__2052;
wire            n594____DOLLAR__2045;
wire            n595____DOLLAR__2038;
wire            n596____DOLLAR__2031;
wire            n597____DOLLAR__2024;
wire            n598____DOLLAR__2017;
wire            n599____DOLLAR__2010;
wire     [39:0] n59____DOLLAR__2925;
wire            n5____DOLLAR__504;
wire            n600____DOLLAR__2003;
wire            n601____DOLLAR__1996;
wire            n602____DOLLAR__1989;
wire            n603____DOLLAR__1982;
wire            n604____DOLLAR__1975;
wire            n605____DOLLAR__1968;
wire            n606____DOLLAR__1961;
wire     [31:0] n607____DOLLAR__1963;
wire     [31:0] n608____DOLLAR__1970;
wire     [31:0] n609____DOLLAR__1977;
wire     [63:0] n60____DOLLAR__2933;
wire     [31:0] n610____DOLLAR__1984;
wire     [31:0] n611____DOLLAR__1991;
wire     [31:0] n612____DOLLAR__1998;
wire     [31:0] n613____DOLLAR__2005;
wire     [31:0] n614____DOLLAR__2012;
wire     [31:0] n615____DOLLAR__2019;
wire     [31:0] n616____DOLLAR__2026;
wire     [31:0] n617____DOLLAR__2033;
wire     [31:0] n618____DOLLAR__2040;
wire     [31:0] n619____DOLLAR__2047;
wire            n61____DOLLAR__3109;
wire     [31:0] n620____DOLLAR__2054;
wire     [31:0] n621____DOLLAR__2061;
wire     [31:0] n622____DOLLAR__1948;
wire     [31:0] n623____DOLLAR__2062;
wire      [7:0] n624____DOLLAR__2071;
wire      [7:0] n625____DOLLAR__2070;
wire      [7:0] n626____DOLLAR__2073;
wire      [7:0] n627____DOLLAR__2074;
wire            n628____DOLLAR__2179;
wire            n629____DOLLAR__2172;
wire     [15:0] n62____DOLLAR__2937;
wire            n630____DOLLAR__2165;
wire            n631____DOLLAR__2158;
wire            n632____DOLLAR__2151;
wire            n633____DOLLAR__2144;
wire            n634____DOLLAR__2137;
wire            n635____DOLLAR__2130;
wire            n636____DOLLAR__2123;
wire            n637____DOLLAR__2116;
wire            n638____DOLLAR__2109;
wire            n639____DOLLAR__2102;
wire     [47:0] n63____DOLLAR__2935;
wire            n640____DOLLAR__2095;
wire            n641____DOLLAR__2088;
wire            n642____DOLLAR__2081;
wire     [31:0] n643____DOLLAR__2083;
wire     [31:0] n644____DOLLAR__2090;
wire     [31:0] n645____DOLLAR__2097;
wire     [31:0] n646____DOLLAR__2104;
wire     [31:0] n647____DOLLAR__2111;
wire     [31:0] n648____DOLLAR__2118;
wire     [31:0] n649____DOLLAR__2125;
wire     [63:0] n64____DOLLAR__2943;
wire     [31:0] n650____DOLLAR__2132;
wire     [31:0] n651____DOLLAR__2139;
wire     [31:0] n652____DOLLAR__2146;
wire     [31:0] n653____DOLLAR__2153;
wire     [31:0] n654____DOLLAR__2160;
wire     [31:0] n655____DOLLAR__2167;
wire     [31:0] n656____DOLLAR__2174;
wire     [31:0] n657____DOLLAR__2181;
wire     [31:0] n658____DOLLAR__2065;
wire     [31:0] n659____DOLLAR__2182;
wire      [7:0] n65____DOLLAR__2947;
wire      [7:0] n660____DOLLAR__2190;
wire      [7:0] n661____DOLLAR__2183;
wire      [7:0] n662____DOLLAR__2192;
wire      [7:0] n663____DOLLAR__2193;
wire            n664____DOLLAR__2298;
wire            n665____DOLLAR__2291;
wire            n666____DOLLAR__2284;
wire            n667____DOLLAR__2277;
wire            n668____DOLLAR__2270;
wire            n669____DOLLAR__2263;
wire     [55:0] n66____DOLLAR__2945;
wire            n670____DOLLAR__2256;
wire            n671____DOLLAR__2249;
wire            n672____DOLLAR__2242;
wire            n673____DOLLAR__2235;
wire            n674____DOLLAR__2228;
wire            n675____DOLLAR__2221;
wire            n676____DOLLAR__2214;
wire            n677____DOLLAR__2207;
wire            n678____DOLLAR__2200;
wire     [31:0] n679____DOLLAR__2202;
wire     [63:0] n67____DOLLAR__2953;
wire     [31:0] n680____DOLLAR__2209;
wire     [31:0] n681____DOLLAR__2216;
wire     [31:0] n682____DOLLAR__2223;
wire     [31:0] n683____DOLLAR__2230;
wire     [31:0] n684____DOLLAR__2237;
wire     [31:0] n685____DOLLAR__2244;
wire     [31:0] n686____DOLLAR__2251;
wire     [31:0] n687____DOLLAR__2258;
wire     [31:0] n688____DOLLAR__2265;
wire     [31:0] n689____DOLLAR__2272;
wire     [63:0] n68____DOLLAR__3111;
wire     [31:0] n690____DOLLAR__2279;
wire     [31:0] n691____DOLLAR__2286;
wire     [31:0] n692____DOLLAR__2293;
wire     [31:0] n693____DOLLAR__2300;
wire     [31:0] n694____DOLLAR__2187;
wire     [31:0] n695____DOLLAR__2301;
wire      [7:0] n696____DOLLAR__2310;
wire      [7:0] n697____DOLLAR__2309;
wire      [7:0] n698____DOLLAR__2312;
wire      [7:0] n699____DOLLAR__2313;
wire     [63:0] n69____DOLLAR__3116;
wire     [12:0] n6____DOLLAR__501;
wire            n700____DOLLAR__2418;
wire            n701____DOLLAR__2411;
wire            n702____DOLLAR__2404;
wire            n703____DOLLAR__2397;
wire            n704____DOLLAR__2390;
wire            n705____DOLLAR__2383;
wire            n706____DOLLAR__2376;
wire            n707____DOLLAR__2369;
wire            n708____DOLLAR__2362;
wire            n709____DOLLAR__2355;
wire     [63:0] n70____DOLLAR__3121;
wire            n710____DOLLAR__2348;
wire            n711____DOLLAR__2341;
wire            n712____DOLLAR__2334;
wire            n713____DOLLAR__2327;
wire            n714____DOLLAR__2320;
wire     [31:0] n715____DOLLAR__2322;
wire     [31:0] n716____DOLLAR__2329;
wire     [31:0] n717____DOLLAR__2336;
wire     [31:0] n718____DOLLAR__2343;
wire     [31:0] n719____DOLLAR__2350;
wire     [63:0] n71____DOLLAR__3126;
wire     [31:0] n720____DOLLAR__2357;
wire     [31:0] n721____DOLLAR__2364;
wire     [31:0] n722____DOLLAR__2371;
wire     [31:0] n723____DOLLAR__2378;
wire     [31:0] n724____DOLLAR__2385;
wire     [31:0] n725____DOLLAR__2392;
wire     [31:0] n726____DOLLAR__2399;
wire     [31:0] n727____DOLLAR__2406;
wire     [31:0] n728____DOLLAR__2413;
wire     [31:0] n729____DOLLAR__2420;
wire     [63:0] n72____DOLLAR__3131;
wire     [31:0] n730____DOLLAR__2304;
wire     [31:0] n731____DOLLAR__2421;
wire      [7:0] n732____DOLLAR__2429;
wire      [7:0] n733____DOLLAR__2422;
wire      [7:0] n734____DOLLAR__2431;
wire      [7:0] n735____DOLLAR__2432;
wire            n736____DOLLAR__2537;
wire            n737____DOLLAR__2530;
wire            n738____DOLLAR__2523;
wire            n739____DOLLAR__2516;
wire     [63:0] n73____DOLLAR__3136;
wire            n740____DOLLAR__2509;
wire            n741____DOLLAR__2502;
wire            n742____DOLLAR__2495;
wire            n743____DOLLAR__2488;
wire            n744____DOLLAR__2481;
wire            n745____DOLLAR__2474;
wire            n746____DOLLAR__2467;
wire            n747____DOLLAR__2460;
wire            n748____DOLLAR__2453;
wire            n749____DOLLAR__2446;
wire     [63:0] n74____DOLLAR__3141;
wire            n750____DOLLAR__2439;
wire     [31:0] n751____DOLLAR__2441;
wire     [31:0] n752____DOLLAR__2448;
wire     [31:0] n753____DOLLAR__2455;
wire     [31:0] n754____DOLLAR__2462;
wire     [31:0] n755____DOLLAR__2469;
wire     [31:0] n756____DOLLAR__2476;
wire     [31:0] n757____DOLLAR__2483;
wire     [31:0] n758____DOLLAR__2490;
wire     [31:0] n759____DOLLAR__2497;
wire            n75____DOLLAR__3104;
wire     [31:0] n760____DOLLAR__2504;
wire     [31:0] n761____DOLLAR__2511;
wire     [31:0] n762____DOLLAR__2518;
wire     [31:0] n763____DOLLAR__2525;
wire     [31:0] n764____DOLLAR__2532;
wire     [31:0] n765____DOLLAR__2539;
wire     [31:0] n766____DOLLAR__2426;
wire     [31:0] n767____DOLLAR__2540;
wire      [7:0] n768____DOLLAR__2549;
wire      [7:0] n769____DOLLAR__2548;
wire            n76____DOLLAR__3099;
wire      [7:0] n770____DOLLAR__2551;
wire      [7:0] n771____DOLLAR__2552;
wire            n772____DOLLAR__2657;
wire            n773____DOLLAR__2650;
wire            n774____DOLLAR__2643;
wire            n775____DOLLAR__2636;
wire            n776____DOLLAR__2629;
wire            n777____DOLLAR__2622;
wire            n778____DOLLAR__2615;
wire            n779____DOLLAR__2608;
wire     [63:0] n77____DOLLAR__2961;
wire            n780____DOLLAR__2601;
wire            n781____DOLLAR__2594;
wire            n782____DOLLAR__2587;
wire            n783____DOLLAR__2580;
wire            n784____DOLLAR__2573;
wire            n785____DOLLAR__2566;
wire            n786____DOLLAR__2559;
wire     [31:0] n787____DOLLAR__2561;
wire     [31:0] n788____DOLLAR__2568;
wire     [31:0] n789____DOLLAR__2575;
wire            n78____DOLLAR__3094;
wire     [31:0] n790____DOLLAR__2582;
wire     [31:0] n791____DOLLAR__2589;
wire     [31:0] n792____DOLLAR__2596;
wire     [31:0] n793____DOLLAR__2603;
wire     [31:0] n794____DOLLAR__2610;
wire     [31:0] n795____DOLLAR__2617;
wire     [31:0] n796____DOLLAR__2624;
wire     [31:0] n797____DOLLAR__2631;
wire     [31:0] n798____DOLLAR__2638;
wire     [31:0] n799____DOLLAR__2645;
wire     [63:0] n79____DOLLAR__2971;
wire     [12:0] n7____DOLLAR__506;
wire     [31:0] n800____DOLLAR__2652;
wire     [31:0] n801____DOLLAR__2659;
wire     [31:0] n802____DOLLAR__2543;
wire     [31:0] n803____DOLLAR__2660;
wire     [31:0] n804____DOLLAR__2665;
wire            n80____DOLLAR__3089;
wire     [63:0] n81____DOLLAR__2981;
wire            n82____DOLLAR__3084;
wire     [63:0] n83____DOLLAR__2991;
wire            n84____DOLLAR__3079;
wire     [63:0] n85____DOLLAR__3001;
wire            n86____DOLLAR__3074;
wire     [55:0] n87____DOLLAR__3013;
wire      [7:0] n88____DOLLAR__3003;
wire     [63:0] n89____DOLLAR__3019;
wire            n8____DOLLAR__496;
wire            n90____DOLLAR__3069;
wire     [47:0] n91____DOLLAR__3031;
wire     [15:0] n92____DOLLAR__3021;
wire     [63:0] n93____DOLLAR__3037;
wire     [39:0] n94____DOLLAR__3049;
wire     [23:0] n95____DOLLAR__3039;
wire     [63:0] n96____DOLLAR__3055;
wire     [63:0] n97____DOLLAR__3071;
wire     [63:0] n98____DOLLAR__3076;
wire     [63:0] n99____DOLLAR__3081;
wire            n9____DOLLAR__491;
wire            rst;
reg     [63:0] TXFIFO_BUFF[31:0];
assign TXFIFO_BUFF_0 = TXFIFO_BUFF[0] ;
assign TXFIFO_BUFF_1 = TXFIFO_BUFF[1] ;
assign TXFIFO_BUFF_2 = TXFIFO_BUFF[2] ;
assign TXFIFO_BUFF_3 = TXFIFO_BUFF[3] ;
assign TXFIFO_BUFF_4 = TXFIFO_BUFF[4] ;
assign TXFIFO_BUFF_5 = TXFIFO_BUFF[5] ;
assign TXFIFO_BUFF_6 = TXFIFO_BUFF[6] ;
assign TXFIFO_BUFF_7 = TXFIFO_BUFF[7] ;
assign TXFIFO_BUFF_8 = TXFIFO_BUFF[8] ;
assign TXFIFO_BUFF_9 = TXFIFO_BUFF[9] ;
assign TXFIFO_BUFF_10 = TXFIFO_BUFF[10] ;
assign TXFIFO_BUFF_11 = TXFIFO_BUFF[11] ;
assign TXFIFO_BUFF_12 = TXFIFO_BUFF[12] ;
assign TXFIFO_BUFF_13 = TXFIFO_BUFF[13] ;
assign TXFIFO_BUFF_14 = TXFIFO_BUFF[14] ;
assign TXFIFO_BUFF_15 = TXFIFO_BUFF[15] ;
assign TXFIFO_BUFF_16 = TXFIFO_BUFF[16] ;
assign TXFIFO_BUFF_17 = TXFIFO_BUFF[17] ;
assign TXFIFO_BUFF_18 = TXFIFO_BUFF[18] ;
assign TXFIFO_BUFF_19 = TXFIFO_BUFF[19] ;
assign TXFIFO_BUFF_20 = TXFIFO_BUFF[20] ;
assign TXFIFO_BUFF_21 = TXFIFO_BUFF[21] ;
assign TXFIFO_BUFF_22 = TXFIFO_BUFF[22] ;
assign TXFIFO_BUFF_23 = TXFIFO_BUFF[23] ;
assign TXFIFO_BUFF_24 = TXFIFO_BUFF[24] ;
assign TXFIFO_BUFF_25 = TXFIFO_BUFF[25] ;
assign TXFIFO_BUFF_26 = TXFIFO_BUFF[26] ;
assign TXFIFO_BUFF_27 = TXFIFO_BUFF[27] ;
assign TXFIFO_BUFF_28 = TXFIFO_BUFF[28] ;
assign TXFIFO_BUFF_29 = TXFIFO_BUFF[29] ;
assign TXFIFO_BUFF_30 = TXFIFO_BUFF[30] ;
assign TXFIFO_BUFF_31 = TXFIFO_BUFF[31] ;
assign n0____DOLLAR__124 =  ( RESETN ) == ( 1'b1 )  ;
assign __ILA_TX_FUNC_valid__ = n0____DOLLAR__124 ;
assign n1____DOLLAR__467 =  ( MODE_10G ) == ( 1'b1 )  ;
assign n2____DOLLAR__472 =  ( TX_STATE ) == ( 5'd8 )  ;
assign n3____DOLLAR__474 =  ( n1____DOLLAR__467 ) & (n2____DOLLAR__472 )  ;
assign __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ = n3____DOLLAR__474 ;
assign n5____DOLLAR__504 =  $signed( TX_WCNT ) > $signed( 16'd0 )  ;
assign n6____DOLLAR__501 =  ( TXFIFO_WUSED_QWD ) - ( 13'd1 )  ;
assign n7____DOLLAR__506 =  ( n5____DOLLAR__504 ) ? ( n6____DOLLAR__501 ) : ( TXFIFO_WUSED_QWD ) ;
assign n8____DOLLAR__496 =  $signed( TX_WCNT ) > $signed( 16'd0 )  ;
assign n9____DOLLAR__491 =  ( TXFIFO_BUFF_RD_PTR ) == ( 5'd16 )  ;
assign n10____DOLLAR__486 =  ( TXFIFO_BUFF_RD_PTR ) + ( 5'd1 )  ;
assign n11____DOLLAR__493 =  ( n9____DOLLAR__491 ) ? ( 5'd0 ) : ( n10____DOLLAR__486 ) ;
assign n12____DOLLAR__498 =  ( n8____DOLLAR__496 ) ? ( n11____DOLLAR__493 ) : ( TXFIFO_BUFF_RD_PTR ) ;
assign n13____DOLLAR__481 =  $signed( TX_WCNT ) > $signed( 16'd0 )  ;
assign n14____DOLLAR__477 =  (  TXFIFO_BUFF [ TXFIFO_BUFF_RD_PTR ] )  ;
assign n15____DOLLAR__483 =  ( n13____DOLLAR__481 ) ? ( n14____DOLLAR__477 ) : ( TXFIFO_RD_OUTPUT ) ;
assign n16____DOLLAR__3169 =  $signed( TX_WCNT ) < $signed( 16'd0 )  ;
assign n17____DOLLAR__3171 =  ( n16____DOLLAR__3169 ) ? ( 5'd8 ) : ( 5'd16 ) ;
assign n18____DOLLAR__3176 =  $signed( TX_WCNT ) < $signed( 16'd16 )  ;
assign n19____DOLLAR__3178 =  ( n18____DOLLAR__3176 ) ? ( 8'd1 ) : ( TX_STATE_ENCAP ) ;
assign n20____DOLLAR__3160 =  ( TX_STATE_ENCAP ) == ( 8'd1 )  ;
assign n21____DOLLAR__3157 =  ( TX_B2B_CNTR ) - ( 6'd1 )  ;
assign n22____DOLLAR__3162 =  ( n20____DOLLAR__3160 ) ? ( n21____DOLLAR__3157 ) : ( TX_B2B_CNTR ) ;
assign n23____DOLLAR__3181 =  ( TX_WCNT ) - ( 16'd8 )  ;
assign n24____DOLLAR__3152 =  $signed( TX_WCNT ) > $signed( 16'd7 )  ;
assign n25____DOLLAR__3144 =  ( TX_WCNT ) == ( 16'd7 )  ;
assign n26____DOLLAR__3146 =  $signed( TX_WCNT ) < $signed( 16'd7 )  ;
assign n27____DOLLAR__3148 =  ( n25____DOLLAR__3144 ) | ( n26____DOLLAR__3146 )  ;
assign n28____DOLLAR__510 = TX_PACKET_BYTE_CNT[2:0] ;
assign n29____DOLLAR__3139 =  ( n28____DOLLAR__510 ) == ( 3'd0 )  ;
assign n30____DOLLAR__3134 =  ( n28____DOLLAR__510 ) == ( 3'd1 )  ;
assign n31____DOLLAR__2739 =  ( $signed( CRC ) >>> ( 32'd24 ))  ;
assign n32____DOLLAR__2740 =  ( n31____DOLLAR__2739 ) & ( 32'd255 )  ;
assign n33____DOLLAR__2733 =  ( $signed( CRC ) >>> ( 32'd8 ))  ;
assign n34____DOLLAR__2734 =  ( n33____DOLLAR__2733 ) & ( 32'd65280 )  ;
assign n35____DOLLAR__2741 =  ( n32____DOLLAR__2740 ) | ( n34____DOLLAR__2734 )  ;
assign n36____DOLLAR__2727 =  ( CRC ) << ( 32'd8 )  ;
assign n37____DOLLAR__2728 =  ( n36____DOLLAR__2727 ) & ( 32'd16711680 )  ;
assign n38____DOLLAR__2742 =  ( n35____DOLLAR__2741 ) | ( n37____DOLLAR__2728 )  ;
assign n39____DOLLAR__2721 =  ( CRC ) << ( 32'd24 )  ;
assign n40____DOLLAR__2717 =  { ( 16'd65280 ) , ( 16'd0 ) }  ;
assign n41____DOLLAR__2722 =  ( n39____DOLLAR__2721 ) & ( n40____DOLLAR__2717 )  ;
assign n42____DOLLAR__2743 =  ( n38____DOLLAR__2742 ) | ( n41____DOLLAR__2722 )  ;
assign n43____DOLLAR__2869 = TXFIFO_RD_OUTPUT[7:0] ;
assign n44____DOLLAR__2875 =  { ( n42____DOLLAR__2743 ) , ( n43____DOLLAR__2869 ) }  ;
assign n45____DOLLAR__2883 =  { ( 24'd460797 ) , ( n44____DOLLAR__2875 ) }  ;
assign n46____DOLLAR__3129 =  ( n28____DOLLAR__510 ) == ( 3'd2 )  ;
assign n47____DOLLAR__2885 = TXFIFO_RD_OUTPUT[15:0] ;
assign n48____DOLLAR__2891 =  { ( n42____DOLLAR__2743 ) , ( n47____DOLLAR__2885 ) }  ;
assign n49____DOLLAR__2899 =  { ( 16'd2045 ) , ( n48____DOLLAR__2891 ) }  ;
assign n50____DOLLAR__3124 =  ( n28____DOLLAR__510 ) == ( 3'd3 )  ;
assign n51____DOLLAR__2901 = TXFIFO_RD_OUTPUT[23:0] ;
assign n52____DOLLAR__2907 =  { ( n42____DOLLAR__2743 ) , ( n51____DOLLAR__2901 ) }  ;
assign n53____DOLLAR__2915 =  { ( 8'd253 ) , ( n52____DOLLAR__2907 ) }  ;
assign n54____DOLLAR__3119 =  ( n28____DOLLAR__510 ) == ( 3'd4 )  ;
assign n55____DOLLAR__2917 = TXFIFO_RD_OUTPUT[31:0] ;
assign n56____DOLLAR__2923 =  { ( n42____DOLLAR__2743 ) , ( n55____DOLLAR__2917 ) }  ;
assign n57____DOLLAR__3114 =  ( n28____DOLLAR__510 ) == ( 3'd5 )  ;
assign n58____DOLLAR__2927 = n42____DOLLAR__2743[23:0] ;
assign n59____DOLLAR__2925 = TXFIFO_RD_OUTPUT[39:0] ;
assign n60____DOLLAR__2933 =  { ( n58____DOLLAR__2927 ) , ( n59____DOLLAR__2925 ) }  ;
assign n61____DOLLAR__3109 =  ( n28____DOLLAR__510 ) == ( 3'd6 )  ;
assign n62____DOLLAR__2937 = n42____DOLLAR__2743[15:0] ;
assign n63____DOLLAR__2935 = TXFIFO_RD_OUTPUT[47:0] ;
assign n64____DOLLAR__2943 =  { ( n62____DOLLAR__2937 ) , ( n63____DOLLAR__2935 ) }  ;
assign n65____DOLLAR__2947 = n42____DOLLAR__2743[7:0] ;
assign n66____DOLLAR__2945 = TXFIFO_RD_OUTPUT[55:0] ;
assign n67____DOLLAR__2953 =  { ( n65____DOLLAR__2947 ) , ( n66____DOLLAR__2945 ) }  ;
assign n68____DOLLAR__3111 =  ( n61____DOLLAR__3109 ) ? ( n64____DOLLAR__2943 ) : ( n67____DOLLAR__2953 ) ;
assign n69____DOLLAR__3116 =  ( n57____DOLLAR__3114 ) ? ( n60____DOLLAR__2933 ) : ( n68____DOLLAR__3111 ) ;
assign n70____DOLLAR__3121 =  ( n54____DOLLAR__3119 ) ? ( n56____DOLLAR__2923 ) : ( n69____DOLLAR__3116 ) ;
assign n71____DOLLAR__3126 =  ( n50____DOLLAR__3124 ) ? ( n53____DOLLAR__2915 ) : ( n70____DOLLAR__3121 ) ;
assign n72____DOLLAR__3131 =  ( n46____DOLLAR__3129 ) ? ( n49____DOLLAR__2899 ) : ( n71____DOLLAR__3126 ) ;
assign n73____DOLLAR__3136 =  ( n30____DOLLAR__3134 ) ? ( n45____DOLLAR__2883 ) : ( n72____DOLLAR__3131 ) ;
assign n74____DOLLAR__3141 =  ( n29____DOLLAR__3139 ) ? ( TXFIFO_RD_OUTPUT ) : ( n73____DOLLAR__3136 ) ;
assign n75____DOLLAR__3104 =  $signed( TX_WCNT ) < $signed( 16'd0 )  ;
assign n76____DOLLAR__3099 =  ( n28____DOLLAR__510 ) == ( 3'd0 )  ;
assign n77____DOLLAR__2961 =  { ( 32'd117901309 ) , ( n42____DOLLAR__2743 ) }  ;
assign n78____DOLLAR__3094 =  ( n28____DOLLAR__510 ) == ( 3'd1 )  ;
assign n79____DOLLAR__2971 =  { ( 32'd117901063 ) , ( 32'd117901063 ) }  ;
assign n80____DOLLAR__3089 =  ( n28____DOLLAR__510 ) == ( 3'd2 )  ;
assign n81____DOLLAR__2981 =  { ( 32'd117901063 ) , ( 32'd117901063 ) }  ;
assign n82____DOLLAR__3084 =  ( n28____DOLLAR__510 ) == ( 3'd3 )  ;
assign n83____DOLLAR__2991 =  { ( 32'd117901063 ) , ( 32'd117901063 ) }  ;
assign n84____DOLLAR__3079 =  ( n28____DOLLAR__510 ) == ( 3'd4 )  ;
assign n85____DOLLAR__3001 =  { ( 32'd117901063 ) , ( 32'd117901309 ) }  ;
assign n86____DOLLAR__3074 =  ( n28____DOLLAR__510 ) == ( 3'd5 )  ;
assign n87____DOLLAR__3013 =  { ( 32'd117901063 ) , ( 24'd460797 ) }  ;
assign n88____DOLLAR__3003 = n42____DOLLAR__2743[31:24] ;
assign n89____DOLLAR__3019 =  { ( n87____DOLLAR__3013 ) , ( n88____DOLLAR__3003 ) }  ;
assign n90____DOLLAR__3069 =  ( n28____DOLLAR__510 ) == ( 3'd6 )  ;
assign n91____DOLLAR__3031 =  { ( 32'd117901063 ) , ( 16'd2045 ) }  ;
assign n92____DOLLAR__3021 = n42____DOLLAR__2743[31:16] ;
assign n93____DOLLAR__3037 =  { ( n91____DOLLAR__3031 ) , ( n92____DOLLAR__3021 ) }  ;
assign n94____DOLLAR__3049 =  { ( 32'd117901063 ) , ( 8'd253 ) }  ;
assign n95____DOLLAR__3039 = n42____DOLLAR__2743[31:8] ;
assign n96____DOLLAR__3055 =  { ( n94____DOLLAR__3049 ) , ( n95____DOLLAR__3039 ) }  ;
assign n97____DOLLAR__3071 =  ( n90____DOLLAR__3069 ) ? ( n93____DOLLAR__3037 ) : ( n96____DOLLAR__3055 ) ;
assign n98____DOLLAR__3076 =  ( n86____DOLLAR__3074 ) ? ( n89____DOLLAR__3019 ) : ( n97____DOLLAR__3071 ) ;
assign n99____DOLLAR__3081 =  ( n84____DOLLAR__3079 ) ? ( n85____DOLLAR__3001 ) : ( n98____DOLLAR__3076 ) ;
assign n100____DOLLAR__3086 =  ( n82____DOLLAR__3084 ) ? ( n83____DOLLAR__2991 ) : ( n99____DOLLAR__3081 ) ;
assign n101____DOLLAR__3091 =  ( n80____DOLLAR__3089 ) ? ( n81____DOLLAR__2981 ) : ( n100____DOLLAR__3086 ) ;
assign n102____DOLLAR__3096 =  ( n78____DOLLAR__3094 ) ? ( n79____DOLLAR__2971 ) : ( n101____DOLLAR__3091 ) ;
assign n103____DOLLAR__3101 =  ( n76____DOLLAR__3099 ) ? ( n77____DOLLAR__2961 ) : ( n102____DOLLAR__3096 ) ;
assign n104____DOLLAR__3065 =  { ( 32'd117901063 ) , ( 32'd117901063 ) }  ;
assign n105____DOLLAR__3106 =  ( n75____DOLLAR__3104 ) ? ( n103____DOLLAR__3101 ) : ( n104____DOLLAR__3065 ) ;
assign n106____DOLLAR__3149 =  ( n27____DOLLAR__3148 ) ? ( n74____DOLLAR__3141 ) : ( n105____DOLLAR__3106 ) ;
assign n107____DOLLAR__3154 =  ( n24____DOLLAR__3152 ) ? ( TXFIFO_RD_OUTPUT ) : ( n106____DOLLAR__3149 ) ;
assign n108____DOLLAR__2865 =  $signed( TX_WCNT ) > $signed( 16'd7 )  ;
assign n109____DOLLAR__2855 =  ( TX_WCNT ) == ( 16'd7 )  ;
assign n110____DOLLAR__2857 =  $signed( TX_WCNT ) < $signed( 16'd7 )  ;
assign n111____DOLLAR__2859 =  ( n109____DOLLAR__2855 ) | ( n110____DOLLAR__2857 )  ;
assign n112____DOLLAR__2850 =  ( n28____DOLLAR__510 ) == ( 3'd0 )  ;
assign n113____DOLLAR__2843 =  ( n28____DOLLAR__510 ) == ( 3'd1 )  ;
assign n114____DOLLAR__2836 =  ( n28____DOLLAR__510 ) == ( 3'd2 )  ;
assign n115____DOLLAR__2829 =  ( n28____DOLLAR__510 ) == ( 3'd3 )  ;
assign n116____DOLLAR__2822 =  ( n28____DOLLAR__510 ) == ( 3'd4 )  ;
assign n117____DOLLAR__2815 =  ( n28____DOLLAR__510 ) == ( 3'd5 )  ;
assign n118____DOLLAR__2808 =  ( n28____DOLLAR__510 ) == ( 3'd6 )  ;
assign n119____DOLLAR__2810 =  ( n118____DOLLAR__2808 ) ? ( 8'd0 ) : ( 8'd0 ) ;
assign n120____DOLLAR__2817 =  ( n117____DOLLAR__2815 ) ? ( 8'd0 ) : ( n119____DOLLAR__2810 ) ;
assign n121____DOLLAR__2824 =  ( n116____DOLLAR__2822 ) ? ( 8'd0 ) : ( n120____DOLLAR__2817 ) ;
assign n122____DOLLAR__2831 =  ( n115____DOLLAR__2829 ) ? ( 8'd128 ) : ( n121____DOLLAR__2824 ) ;
assign n123____DOLLAR__2838 =  ( n114____DOLLAR__2836 ) ? ( 8'd192 ) : ( n122____DOLLAR__2831 ) ;
assign n124____DOLLAR__2845 =  ( n113____DOLLAR__2843 ) ? ( 8'd224 ) : ( n123____DOLLAR__2838 ) ;
assign n125____DOLLAR__2852 =  ( n112____DOLLAR__2850 ) ? ( 8'd0 ) : ( n124____DOLLAR__2845 ) ;
assign n126____DOLLAR__2799 =  $signed( TX_WCNT ) < $signed( 16'd0 )  ;
assign n127____DOLLAR__2794 =  ( n28____DOLLAR__510 ) == ( 3'd0 )  ;
assign n128____DOLLAR__2787 =  ( n28____DOLLAR__510 ) == ( 3'd1 )  ;
assign n129____DOLLAR__2780 =  ( n28____DOLLAR__510 ) == ( 3'd2 )  ;
assign n130____DOLLAR__2773 =  ( n28____DOLLAR__510 ) == ( 3'd3 )  ;
assign n131____DOLLAR__2766 =  ( n28____DOLLAR__510 ) == ( 3'd4 )  ;
assign n132____DOLLAR__2759 =  ( n28____DOLLAR__510 ) == ( 3'd5 )  ;
assign n133____DOLLAR__2752 =  ( n28____DOLLAR__510 ) == ( 3'd6 )  ;
assign n134____DOLLAR__2754 =  ( n133____DOLLAR__2752 ) ? ( 8'd252 ) : ( 8'd248 ) ;
assign n135____DOLLAR__2761 =  ( n132____DOLLAR__2759 ) ? ( 8'd254 ) : ( n134____DOLLAR__2754 ) ;
assign n136____DOLLAR__2768 =  ( n131____DOLLAR__2766 ) ? ( 8'd255 ) : ( n135____DOLLAR__2761 ) ;
assign n137____DOLLAR__2775 =  ( n130____DOLLAR__2773 ) ? ( 8'd255 ) : ( n136____DOLLAR__2768 ) ;
assign n138____DOLLAR__2782 =  ( n129____DOLLAR__2780 ) ? ( 8'd255 ) : ( n137____DOLLAR__2775 ) ;
assign n139____DOLLAR__2789 =  ( n128____DOLLAR__2787 ) ? ( 8'd255 ) : ( n138____DOLLAR__2782 ) ;
assign n140____DOLLAR__2796 =  ( n127____DOLLAR__2794 ) ? ( 8'd240 ) : ( n139____DOLLAR__2789 ) ;
assign n141____DOLLAR__2801 =  ( n126____DOLLAR__2799 ) ? ( n140____DOLLAR__2796 ) : ( 8'd255 ) ;
assign n142____DOLLAR__2860 =  ( n111____DOLLAR__2859 ) ? ( n125____DOLLAR__2852 ) : ( n141____DOLLAR__2801 ) ;
assign n143____DOLLAR__2867 =  ( n108____DOLLAR__2865 ) ? ( 8'd0 ) : ( n142____DOLLAR__2860 ) ;
assign n144____DOLLAR__2705 =  $signed( TX_WCNT ) > $signed( 16'd0 )  ;
assign n145____DOLLAR__2696 =  ( $signed( CRC_IN ) >>> ( 32'd24 ))  ;
assign n146____DOLLAR__2697 =  ( n145____DOLLAR__2696 ) & ( 32'd255 )  ;
assign n147____DOLLAR__2690 =  ( $signed( CRC_IN ) >>> ( 32'd8 ))  ;
assign n148____DOLLAR__2691 =  ( n147____DOLLAR__2690 ) & ( 32'd65280 )  ;
assign n149____DOLLAR__2698 =  ( n146____DOLLAR__2697 ) | ( n148____DOLLAR__2691 )  ;
assign n150____DOLLAR__2684 =  ( CRC_IN ) << ( 32'd8 )  ;
assign n151____DOLLAR__2685 =  ( n150____DOLLAR__2684 ) & ( 32'd16711680 )  ;
assign n152____DOLLAR__2699 =  ( n149____DOLLAR__2698 ) | ( n151____DOLLAR__2685 )  ;
assign n153____DOLLAR__2678 =  ( CRC_IN ) << ( 32'd24 )  ;
assign n154____DOLLAR__2674 =  { ( 16'd65280 ) , ( 16'd0 ) }  ;
assign n155____DOLLAR__2679 =  ( n153____DOLLAR__2678 ) & ( n154____DOLLAR__2674 )  ;
assign n156____DOLLAR__2700 =  ( n152____DOLLAR__2699 ) | ( n155____DOLLAR__2679 )  ;
assign n157____DOLLAR__2701 = ~ ( n156____DOLLAR__2700 ) ;
assign n158____DOLLAR__2707 =  ( n144____DOLLAR__2705 ) ? ( n157____DOLLAR__2701 ) : ( CRC ) ;
assign n159____DOLLAR__508 =  ( TX_WCNT ) == ( TX_WCNT_INI )  ;
assign n160____DOLLAR__743 =  ( n28____DOLLAR__510 ) == ( 3'd0 )  ;
assign n161____DOLLAR__738 =  ( n28____DOLLAR__510 ) == ( 3'd1 )  ;
assign n162____DOLLAR__728 = TXFIFO_RD_OUTPUT[7:0] ;
assign n163____DOLLAR__726 =  { ( 32'd0 ) , ( 24'd0 ) }  ;
assign n164____DOLLAR__734 =  { ( n162____DOLLAR__728 ) , ( n163____DOLLAR__726 ) }  ;
assign n165____DOLLAR__715 =  ( n28____DOLLAR__510 ) == ( 3'd2 )  ;
assign n166____DOLLAR__705 = TXFIFO_RD_OUTPUT[15:0] ;
assign n167____DOLLAR__703 =  { ( 32'd0 ) , ( 16'd0 ) }  ;
assign n168____DOLLAR__711 =  { ( n166____DOLLAR__705 ) , ( n167____DOLLAR__703 ) }  ;
assign n169____DOLLAR__692 =  ( n28____DOLLAR__510 ) == ( 3'd3 )  ;
assign n170____DOLLAR__682 = TXFIFO_RD_OUTPUT[23:0] ;
assign n171____DOLLAR__680 =  { ( 32'd0 ) , ( 8'd0 ) }  ;
assign n172____DOLLAR__688 =  { ( n170____DOLLAR__682 ) , ( n171____DOLLAR__680 ) }  ;
assign n173____DOLLAR__669 =  ( n28____DOLLAR__510 ) == ( 3'd4 )  ;
assign n174____DOLLAR__659 = TXFIFO_RD_OUTPUT[31:0] ;
assign n175____DOLLAR__665 =  { ( n174____DOLLAR__659 ) , ( 32'd0 ) }  ;
assign n176____DOLLAR__654 =  ( n28____DOLLAR__510 ) == ( 3'd5 )  ;
assign n177____DOLLAR__644 = TXFIFO_RD_OUTPUT[39:0] ;
assign n178____DOLLAR__650 =  { ( n177____DOLLAR__644 ) , ( 24'd0 ) }  ;
assign n179____DOLLAR__639 =  ( n28____DOLLAR__510 ) == ( 3'd6 )  ;
assign n180____DOLLAR__629 = TXFIFO_RD_OUTPUT[47:0] ;
assign n181____DOLLAR__635 =  { ( n180____DOLLAR__629 ) , ( 16'd0 ) }  ;
assign n182____DOLLAR__619 = TXFIFO_RD_OUTPUT[55:0] ;
assign n183____DOLLAR__625 =  { ( n182____DOLLAR__619 ) , ( 8'd0 ) }  ;
assign n184____DOLLAR__641 =  ( n179____DOLLAR__639 ) ? ( n181____DOLLAR__635 ) : ( n183____DOLLAR__625 ) ;
assign n185____DOLLAR__656 =  ( n176____DOLLAR__654 ) ? ( n178____DOLLAR__650 ) : ( n184____DOLLAR__641 ) ;
assign n186____DOLLAR__671 =  ( n173____DOLLAR__669 ) ? ( n175____DOLLAR__665 ) : ( n185____DOLLAR__656 ) ;
assign n187____DOLLAR__694 =  ( n169____DOLLAR__692 ) ? ( n172____DOLLAR__688 ) : ( n186____DOLLAR__671 ) ;
assign n188____DOLLAR__717 =  ( n165____DOLLAR__715 ) ? ( n168____DOLLAR__711 ) : ( n187____DOLLAR__694 ) ;
assign n189____DOLLAR__740 =  ( n161____DOLLAR__738 ) ? ( n164____DOLLAR__734 ) : ( n188____DOLLAR__717 ) ;
assign n190____DOLLAR__745 =  ( n160____DOLLAR__743 ) ? ( TXFIFO_RD_OUTPUT ) : ( n189____DOLLAR__740 ) ;
assign n191____DOLLAR__614 =  ( n28____DOLLAR__510 ) == ( 3'd0 )  ;
assign n192____DOLLAR__609 =  ( n28____DOLLAR__510 ) == ( 3'd1 )  ;
assign n193____DOLLAR__599 = TXFIFO_RD_OUTPUT[7:0] ;
assign n194____DOLLAR__597 = TX_BUF[63:8] ;
assign n195____DOLLAR__605 =  { ( n193____DOLLAR__599 ) , ( n194____DOLLAR__597 ) }  ;
assign n196____DOLLAR__594 =  ( n28____DOLLAR__510 ) == ( 3'd2 )  ;
assign n197____DOLLAR__584 = TXFIFO_RD_OUTPUT[15:0] ;
assign n198____DOLLAR__582 = TX_BUF[63:16] ;
assign n199____DOLLAR__590 =  { ( n197____DOLLAR__584 ) , ( n198____DOLLAR__582 ) }  ;
assign n200____DOLLAR__579 =  ( n28____DOLLAR__510 ) == ( 3'd3 )  ;
assign n201____DOLLAR__569 = TXFIFO_RD_OUTPUT[23:0] ;
assign n202____DOLLAR__567 = TX_BUF[63:24] ;
assign n203____DOLLAR__575 =  { ( n201____DOLLAR__569 ) , ( n202____DOLLAR__567 ) }  ;
assign n204____DOLLAR__564 =  ( n28____DOLLAR__510 ) == ( 3'd4 )  ;
assign n205____DOLLAR__554 = TXFIFO_RD_OUTPUT[31:0] ;
assign n206____DOLLAR__552 = TX_BUF[63:32] ;
assign n207____DOLLAR__560 =  { ( n205____DOLLAR__554 ) , ( n206____DOLLAR__552 ) }  ;
assign n208____DOLLAR__549 =  ( n28____DOLLAR__510 ) == ( 3'd5 )  ;
assign n209____DOLLAR__539 = TXFIFO_RD_OUTPUT[39:0] ;
assign n210____DOLLAR__537 = TX_BUF[63:40] ;
assign n211____DOLLAR__545 =  { ( n209____DOLLAR__539 ) , ( n210____DOLLAR__537 ) }  ;
assign n212____DOLLAR__534 =  ( n28____DOLLAR__510 ) == ( 3'd6 )  ;
assign n213____DOLLAR__524 = TXFIFO_RD_OUTPUT[47:0] ;
assign n214____DOLLAR__522 = TX_BUF[63:48] ;
assign n215____DOLLAR__530 =  { ( n213____DOLLAR__524 ) , ( n214____DOLLAR__522 ) }  ;
assign n216____DOLLAR__514 = TXFIFO_RD_OUTPUT[55:0] ;
assign n217____DOLLAR__512 = TX_BUF[63:56] ;
assign n218____DOLLAR__520 =  { ( n216____DOLLAR__514 ) , ( n217____DOLLAR__512 ) }  ;
assign n219____DOLLAR__536 =  ( n212____DOLLAR__534 ) ? ( n215____DOLLAR__530 ) : ( n218____DOLLAR__520 ) ;
assign n220____DOLLAR__551 =  ( n208____DOLLAR__549 ) ? ( n211____DOLLAR__545 ) : ( n219____DOLLAR__536 ) ;
assign n221____DOLLAR__566 =  ( n204____DOLLAR__564 ) ? ( n207____DOLLAR__560 ) : ( n220____DOLLAR__551 ) ;
assign n222____DOLLAR__581 =  ( n200____DOLLAR__579 ) ? ( n203____DOLLAR__575 ) : ( n221____DOLLAR__566 ) ;
assign n223____DOLLAR__596 =  ( n196____DOLLAR__594 ) ? ( n199____DOLLAR__590 ) : ( n222____DOLLAR__581 ) ;
assign n224____DOLLAR__611 =  ( n192____DOLLAR__609 ) ? ( n195____DOLLAR__605 ) : ( n223____DOLLAR__596 ) ;
assign n225____DOLLAR__616 =  ( n191____DOLLAR__614 ) ? ( TXFIFO_RD_OUTPUT ) : ( n224____DOLLAR__611 ) ;
assign n226____DOLLAR__746 =  ( n159____DOLLAR__508 ) ? ( n190____DOLLAR__745 ) : ( n225____DOLLAR__616 ) ;
assign n227____DOLLAR__2663 =  $signed( TX_WCNT ) > $signed( 16'd0 )  ;
assign n228____DOLLAR__756 = CRC_IN[7:0] ;
assign n229____DOLLAR__749 = CRC_DAT_IN[7:0] ;
assign n230____DOLLAR__758 =  ( n228____DOLLAR__756 ) ^ ( n229____DOLLAR__749 )  ;
assign n231____DOLLAR__759 =  ( n230____DOLLAR__758 ) & ( 8'd15 )  ;
assign n232____DOLLAR__864 =  ( n231____DOLLAR__759 ) == ( 8'd15 )  ;
assign n233____DOLLAR__857 =  ( n231____DOLLAR__759 ) == ( 8'd14 )  ;
assign n234____DOLLAR__850 =  ( n231____DOLLAR__759 ) == ( 8'd13 )  ;
assign n235____DOLLAR__843 =  ( n231____DOLLAR__759 ) == ( 8'd12 )  ;
assign n236____DOLLAR__836 =  ( n231____DOLLAR__759 ) == ( 8'd11 )  ;
assign n237____DOLLAR__829 =  ( n231____DOLLAR__759 ) == ( 8'd10 )  ;
assign n238____DOLLAR__822 =  ( n231____DOLLAR__759 ) == ( 8'd9 )  ;
assign n239____DOLLAR__815 =  ( n231____DOLLAR__759 ) == ( 8'd8 )  ;
assign n240____DOLLAR__808 =  ( n231____DOLLAR__759 ) == ( 8'd7 )  ;
assign n241____DOLLAR__801 =  ( n231____DOLLAR__759 ) == ( 8'd6 )  ;
assign n242____DOLLAR__794 =  ( n231____DOLLAR__759 ) == ( 8'd5 )  ;
assign n243____DOLLAR__787 =  ( n231____DOLLAR__759 ) == ( 8'd4 )  ;
assign n244____DOLLAR__780 =  ( n231____DOLLAR__759 ) == ( 8'd3 )  ;
assign n245____DOLLAR__773 =  ( n231____DOLLAR__759 ) == ( 8'd2 )  ;
assign n246____DOLLAR__766 =  ( n231____DOLLAR__759 ) == ( 8'd1 )  ;
assign n247____DOLLAR__768 =  ( n246____DOLLAR__766 ) ? ( 32'd498536548 ) : ( 32'd0 ) ;
assign n248____DOLLAR__775 =  ( n245____DOLLAR__773 ) ? ( 32'd997073096 ) : ( n247____DOLLAR__768 ) ;
assign n249____DOLLAR__782 =  ( n244____DOLLAR__780 ) ? ( 32'd651767980 ) : ( n248____DOLLAR__775 ) ;
assign n250____DOLLAR__789 =  ( n243____DOLLAR__787 ) ? ( 32'd1994146192 ) : ( n249____DOLLAR__782 ) ;
assign n251____DOLLAR__796 =  ( n242____DOLLAR__794 ) ? ( 32'd1802195444 ) : ( n250____DOLLAR__789 ) ;
assign n252____DOLLAR__803 =  ( n241____DOLLAR__801 ) ? ( 32'd1303535960 ) : ( n251____DOLLAR__796 ) ;
assign n253____DOLLAR__810 =  ( n240____DOLLAR__808 ) ? ( 32'd1342533948 ) : ( n252____DOLLAR__803 ) ;
assign n254____DOLLAR__817 =  ( n239____DOLLAR__815 ) ? ( 32'd-306674912 ) : ( n253____DOLLAR__810 ) ;
assign n255____DOLLAR__824 =  ( n238____DOLLAR__822 ) ? ( 32'd-267414716 ) : ( n254____DOLLAR__817 ) ;
assign n256____DOLLAR__831 =  ( n237____DOLLAR__829 ) ? ( 32'd-690576408 ) : ( n255____DOLLAR__824 ) ;
assign n257____DOLLAR__838 =  ( n236____DOLLAR__836 ) ? ( 32'd-882789492 ) : ( n256____DOLLAR__831 ) ;
assign n258____DOLLAR__845 =  ( n235____DOLLAR__843 ) ? ( 32'd-1687895376 ) : ( n257____DOLLAR__838 ) ;
assign n259____DOLLAR__852 =  ( n234____DOLLAR__850 ) ? ( 32'd-2032938284 ) : ( n258____DOLLAR__845 ) ;
assign n260____DOLLAR__859 =  ( n233____DOLLAR__857 ) ? ( 32'd-1609899400 ) : ( n259____DOLLAR__852 ) ;
assign n261____DOLLAR__866 =  ( n232____DOLLAR__864 ) ? ( 32'd-1111625188 ) : ( n260____DOLLAR__859 ) ;
assign n262____DOLLAR__753 =  ( $signed( CRC_IN ) >>> ( 32'd4 ))  ;
assign n263____DOLLAR__867 =  ( n261____DOLLAR__866 ) ^ ( n262____DOLLAR__753 )  ;
assign n264____DOLLAR__876 = n263____DOLLAR__867[7:0] ;
assign n265____DOLLAR__875 =  ( $signed( n229____DOLLAR__749 ) >>> ( 8'd4 ))  ;
assign n266____DOLLAR__878 =  ( n264____DOLLAR__876 ) ^ ( n265____DOLLAR__875 )  ;
assign n267____DOLLAR__879 =  ( n266____DOLLAR__878 ) & ( 8'd15 )  ;
assign n268____DOLLAR__984 =  ( n267____DOLLAR__879 ) == ( 8'd15 )  ;
assign n269____DOLLAR__977 =  ( n267____DOLLAR__879 ) == ( 8'd14 )  ;
assign n270____DOLLAR__970 =  ( n267____DOLLAR__879 ) == ( 8'd13 )  ;
assign n271____DOLLAR__963 =  ( n267____DOLLAR__879 ) == ( 8'd12 )  ;
assign n272____DOLLAR__956 =  ( n267____DOLLAR__879 ) == ( 8'd11 )  ;
assign n273____DOLLAR__949 =  ( n267____DOLLAR__879 ) == ( 8'd10 )  ;
assign n274____DOLLAR__942 =  ( n267____DOLLAR__879 ) == ( 8'd9 )  ;
assign n275____DOLLAR__935 =  ( n267____DOLLAR__879 ) == ( 8'd8 )  ;
assign n276____DOLLAR__928 =  ( n267____DOLLAR__879 ) == ( 8'd7 )  ;
assign n277____DOLLAR__921 =  ( n267____DOLLAR__879 ) == ( 8'd6 )  ;
assign n278____DOLLAR__914 =  ( n267____DOLLAR__879 ) == ( 8'd5 )  ;
assign n279____DOLLAR__907 =  ( n267____DOLLAR__879 ) == ( 8'd4 )  ;
assign n280____DOLLAR__900 =  ( n267____DOLLAR__879 ) == ( 8'd3 )  ;
assign n281____DOLLAR__893 =  ( n267____DOLLAR__879 ) == ( 8'd2 )  ;
assign n282____DOLLAR__886 =  ( n267____DOLLAR__879 ) == ( 8'd1 )  ;
assign n283____DOLLAR__888 =  ( n282____DOLLAR__886 ) ? ( 32'd498536548 ) : ( 32'd0 ) ;
assign n284____DOLLAR__895 =  ( n281____DOLLAR__893 ) ? ( 32'd997073096 ) : ( n283____DOLLAR__888 ) ;
assign n285____DOLLAR__902 =  ( n280____DOLLAR__900 ) ? ( 32'd651767980 ) : ( n284____DOLLAR__895 ) ;
assign n286____DOLLAR__909 =  ( n279____DOLLAR__907 ) ? ( 32'd1994146192 ) : ( n285____DOLLAR__902 ) ;
assign n287____DOLLAR__916 =  ( n278____DOLLAR__914 ) ? ( 32'd1802195444 ) : ( n286____DOLLAR__909 ) ;
assign n288____DOLLAR__923 =  ( n277____DOLLAR__921 ) ? ( 32'd1303535960 ) : ( n287____DOLLAR__916 ) ;
assign n289____DOLLAR__930 =  ( n276____DOLLAR__928 ) ? ( 32'd1342533948 ) : ( n288____DOLLAR__923 ) ;
assign n290____DOLLAR__937 =  ( n275____DOLLAR__935 ) ? ( 32'd-306674912 ) : ( n289____DOLLAR__930 ) ;
assign n291____DOLLAR__944 =  ( n274____DOLLAR__942 ) ? ( 32'd-267414716 ) : ( n290____DOLLAR__937 ) ;
assign n292____DOLLAR__951 =  ( n273____DOLLAR__949 ) ? ( 32'd-690576408 ) : ( n291____DOLLAR__944 ) ;
assign n293____DOLLAR__958 =  ( n272____DOLLAR__956 ) ? ( 32'd-882789492 ) : ( n292____DOLLAR__951 ) ;
assign n294____DOLLAR__965 =  ( n271____DOLLAR__963 ) ? ( 32'd-1687895376 ) : ( n293____DOLLAR__958 ) ;
assign n295____DOLLAR__972 =  ( n270____DOLLAR__970 ) ? ( 32'd-2032938284 ) : ( n294____DOLLAR__965 ) ;
assign n296____DOLLAR__979 =  ( n269____DOLLAR__977 ) ? ( 32'd-1609899400 ) : ( n295____DOLLAR__972 ) ;
assign n297____DOLLAR__986 =  ( n268____DOLLAR__984 ) ? ( 32'd-1111625188 ) : ( n296____DOLLAR__979 ) ;
assign n298____DOLLAR__870 =  ( $signed( n263____DOLLAR__867 ) >>> ( 32'd4 ))  ;
assign n299____DOLLAR__987 =  ( n297____DOLLAR__986 ) ^ ( n298____DOLLAR__870 )  ;
assign n300____DOLLAR__995 = n299____DOLLAR__987[7:0] ;
assign n301____DOLLAR__988 = CRC_DAT_IN[15:8] ;
assign n302____DOLLAR__997 =  ( n300____DOLLAR__995 ) ^ ( n301____DOLLAR__988 )  ;
assign n303____DOLLAR__998 =  ( n302____DOLLAR__997 ) & ( 8'd15 )  ;
assign n304____DOLLAR__1103 =  ( n303____DOLLAR__998 ) == ( 8'd15 )  ;
assign n305____DOLLAR__1096 =  ( n303____DOLLAR__998 ) == ( 8'd14 )  ;
assign n306____DOLLAR__1089 =  ( n303____DOLLAR__998 ) == ( 8'd13 )  ;
assign n307____DOLLAR__1082 =  ( n303____DOLLAR__998 ) == ( 8'd12 )  ;
assign n308____DOLLAR__1075 =  ( n303____DOLLAR__998 ) == ( 8'd11 )  ;
assign n309____DOLLAR__1068 =  ( n303____DOLLAR__998 ) == ( 8'd10 )  ;
assign n310____DOLLAR__1061 =  ( n303____DOLLAR__998 ) == ( 8'd9 )  ;
assign n311____DOLLAR__1054 =  ( n303____DOLLAR__998 ) == ( 8'd8 )  ;
assign n312____DOLLAR__1047 =  ( n303____DOLLAR__998 ) == ( 8'd7 )  ;
assign n313____DOLLAR__1040 =  ( n303____DOLLAR__998 ) == ( 8'd6 )  ;
assign n314____DOLLAR__1033 =  ( n303____DOLLAR__998 ) == ( 8'd5 )  ;
assign n315____DOLLAR__1026 =  ( n303____DOLLAR__998 ) == ( 8'd4 )  ;
assign n316____DOLLAR__1019 =  ( n303____DOLLAR__998 ) == ( 8'd3 )  ;
assign n317____DOLLAR__1012 =  ( n303____DOLLAR__998 ) == ( 8'd2 )  ;
assign n318____DOLLAR__1005 =  ( n303____DOLLAR__998 ) == ( 8'd1 )  ;
assign n319____DOLLAR__1007 =  ( n318____DOLLAR__1005 ) ? ( 32'd498536548 ) : ( 32'd0 ) ;
assign n320____DOLLAR__1014 =  ( n317____DOLLAR__1012 ) ? ( 32'd997073096 ) : ( n319____DOLLAR__1007 ) ;
assign n321____DOLLAR__1021 =  ( n316____DOLLAR__1019 ) ? ( 32'd651767980 ) : ( n320____DOLLAR__1014 ) ;
assign n322____DOLLAR__1028 =  ( n315____DOLLAR__1026 ) ? ( 32'd1994146192 ) : ( n321____DOLLAR__1021 ) ;
assign n323____DOLLAR__1035 =  ( n314____DOLLAR__1033 ) ? ( 32'd1802195444 ) : ( n322____DOLLAR__1028 ) ;
assign n324____DOLLAR__1042 =  ( n313____DOLLAR__1040 ) ? ( 32'd1303535960 ) : ( n323____DOLLAR__1035 ) ;
assign n325____DOLLAR__1049 =  ( n312____DOLLAR__1047 ) ? ( 32'd1342533948 ) : ( n324____DOLLAR__1042 ) ;
assign n326____DOLLAR__1056 =  ( n311____DOLLAR__1054 ) ? ( 32'd-306674912 ) : ( n325____DOLLAR__1049 ) ;
assign n327____DOLLAR__1063 =  ( n310____DOLLAR__1061 ) ? ( 32'd-267414716 ) : ( n326____DOLLAR__1056 ) ;
assign n328____DOLLAR__1070 =  ( n309____DOLLAR__1068 ) ? ( 32'd-690576408 ) : ( n327____DOLLAR__1063 ) ;
assign n329____DOLLAR__1077 =  ( n308____DOLLAR__1075 ) ? ( 32'd-882789492 ) : ( n328____DOLLAR__1070 ) ;
assign n330____DOLLAR__1084 =  ( n307____DOLLAR__1082 ) ? ( 32'd-1687895376 ) : ( n329____DOLLAR__1077 ) ;
assign n331____DOLLAR__1091 =  ( n306____DOLLAR__1089 ) ? ( 32'd-2032938284 ) : ( n330____DOLLAR__1084 ) ;
assign n332____DOLLAR__1098 =  ( n305____DOLLAR__1096 ) ? ( 32'd-1609899400 ) : ( n331____DOLLAR__1091 ) ;
assign n333____DOLLAR__1105 =  ( n304____DOLLAR__1103 ) ? ( 32'd-1111625188 ) : ( n332____DOLLAR__1098 ) ;
assign n334____DOLLAR__992 =  ( $signed( n299____DOLLAR__987 ) >>> ( 32'd4 ))  ;
assign n335____DOLLAR__1106 =  ( n333____DOLLAR__1105 ) ^ ( n334____DOLLAR__992 )  ;
assign n336____DOLLAR__1115 = n335____DOLLAR__1106[7:0] ;
assign n337____DOLLAR__1114 =  ( $signed( n301____DOLLAR__988 ) >>> ( 8'd4 ))  ;
assign n338____DOLLAR__1117 =  ( n336____DOLLAR__1115 ) ^ ( n337____DOLLAR__1114 )  ;
assign n339____DOLLAR__1118 =  ( n338____DOLLAR__1117 ) & ( 8'd15 )  ;
assign n340____DOLLAR__1223 =  ( n339____DOLLAR__1118 ) == ( 8'd15 )  ;
assign n341____DOLLAR__1216 =  ( n339____DOLLAR__1118 ) == ( 8'd14 )  ;
assign n342____DOLLAR__1209 =  ( n339____DOLLAR__1118 ) == ( 8'd13 )  ;
assign n343____DOLLAR__1202 =  ( n339____DOLLAR__1118 ) == ( 8'd12 )  ;
assign n344____DOLLAR__1195 =  ( n339____DOLLAR__1118 ) == ( 8'd11 )  ;
assign n345____DOLLAR__1188 =  ( n339____DOLLAR__1118 ) == ( 8'd10 )  ;
assign n346____DOLLAR__1181 =  ( n339____DOLLAR__1118 ) == ( 8'd9 )  ;
assign n347____DOLLAR__1174 =  ( n339____DOLLAR__1118 ) == ( 8'd8 )  ;
assign n348____DOLLAR__1167 =  ( n339____DOLLAR__1118 ) == ( 8'd7 )  ;
assign n349____DOLLAR__1160 =  ( n339____DOLLAR__1118 ) == ( 8'd6 )  ;
assign n350____DOLLAR__1153 =  ( n339____DOLLAR__1118 ) == ( 8'd5 )  ;
assign n351____DOLLAR__1146 =  ( n339____DOLLAR__1118 ) == ( 8'd4 )  ;
assign n352____DOLLAR__1139 =  ( n339____DOLLAR__1118 ) == ( 8'd3 )  ;
assign n353____DOLLAR__1132 =  ( n339____DOLLAR__1118 ) == ( 8'd2 )  ;
assign n354____DOLLAR__1125 =  ( n339____DOLLAR__1118 ) == ( 8'd1 )  ;
assign n355____DOLLAR__1127 =  ( n354____DOLLAR__1125 ) ? ( 32'd498536548 ) : ( 32'd0 ) ;
assign n356____DOLLAR__1134 =  ( n353____DOLLAR__1132 ) ? ( 32'd997073096 ) : ( n355____DOLLAR__1127 ) ;
assign n357____DOLLAR__1141 =  ( n352____DOLLAR__1139 ) ? ( 32'd651767980 ) : ( n356____DOLLAR__1134 ) ;
assign n358____DOLLAR__1148 =  ( n351____DOLLAR__1146 ) ? ( 32'd1994146192 ) : ( n357____DOLLAR__1141 ) ;
assign n359____DOLLAR__1155 =  ( n350____DOLLAR__1153 ) ? ( 32'd1802195444 ) : ( n358____DOLLAR__1148 ) ;
assign n360____DOLLAR__1162 =  ( n349____DOLLAR__1160 ) ? ( 32'd1303535960 ) : ( n359____DOLLAR__1155 ) ;
assign n361____DOLLAR__1169 =  ( n348____DOLLAR__1167 ) ? ( 32'd1342533948 ) : ( n360____DOLLAR__1162 ) ;
assign n362____DOLLAR__1176 =  ( n347____DOLLAR__1174 ) ? ( 32'd-306674912 ) : ( n361____DOLLAR__1169 ) ;
assign n363____DOLLAR__1183 =  ( n346____DOLLAR__1181 ) ? ( 32'd-267414716 ) : ( n362____DOLLAR__1176 ) ;
assign n364____DOLLAR__1190 =  ( n345____DOLLAR__1188 ) ? ( 32'd-690576408 ) : ( n363____DOLLAR__1183 ) ;
assign n365____DOLLAR__1197 =  ( n344____DOLLAR__1195 ) ? ( 32'd-882789492 ) : ( n364____DOLLAR__1190 ) ;
assign n366____DOLLAR__1204 =  ( n343____DOLLAR__1202 ) ? ( 32'd-1687895376 ) : ( n365____DOLLAR__1197 ) ;
assign n367____DOLLAR__1211 =  ( n342____DOLLAR__1209 ) ? ( 32'd-2032938284 ) : ( n366____DOLLAR__1204 ) ;
assign n368____DOLLAR__1218 =  ( n341____DOLLAR__1216 ) ? ( 32'd-1609899400 ) : ( n367____DOLLAR__1211 ) ;
assign n369____DOLLAR__1225 =  ( n340____DOLLAR__1223 ) ? ( 32'd-1111625188 ) : ( n368____DOLLAR__1218 ) ;
assign n370____DOLLAR__1109 =  ( $signed( n335____DOLLAR__1106 ) >>> ( 32'd4 ))  ;
assign n371____DOLLAR__1226 =  ( n369____DOLLAR__1225 ) ^ ( n370____DOLLAR__1109 )  ;
assign n372____DOLLAR__1234 = n371____DOLLAR__1226[7:0] ;
assign n373____DOLLAR__1227 = CRC_DAT_IN[23:16] ;
assign n374____DOLLAR__1236 =  ( n372____DOLLAR__1234 ) ^ ( n373____DOLLAR__1227 )  ;
assign n375____DOLLAR__1237 =  ( n374____DOLLAR__1236 ) & ( 8'd15 )  ;
assign n376____DOLLAR__1342 =  ( n375____DOLLAR__1237 ) == ( 8'd15 )  ;
assign n377____DOLLAR__1335 =  ( n375____DOLLAR__1237 ) == ( 8'd14 )  ;
assign n378____DOLLAR__1328 =  ( n375____DOLLAR__1237 ) == ( 8'd13 )  ;
assign n379____DOLLAR__1321 =  ( n375____DOLLAR__1237 ) == ( 8'd12 )  ;
assign n380____DOLLAR__1314 =  ( n375____DOLLAR__1237 ) == ( 8'd11 )  ;
assign n381____DOLLAR__1307 =  ( n375____DOLLAR__1237 ) == ( 8'd10 )  ;
assign n382____DOLLAR__1300 =  ( n375____DOLLAR__1237 ) == ( 8'd9 )  ;
assign n383____DOLLAR__1293 =  ( n375____DOLLAR__1237 ) == ( 8'd8 )  ;
assign n384____DOLLAR__1286 =  ( n375____DOLLAR__1237 ) == ( 8'd7 )  ;
assign n385____DOLLAR__1279 =  ( n375____DOLLAR__1237 ) == ( 8'd6 )  ;
assign n386____DOLLAR__1272 =  ( n375____DOLLAR__1237 ) == ( 8'd5 )  ;
assign n387____DOLLAR__1265 =  ( n375____DOLLAR__1237 ) == ( 8'd4 )  ;
assign n388____DOLLAR__1258 =  ( n375____DOLLAR__1237 ) == ( 8'd3 )  ;
assign n389____DOLLAR__1251 =  ( n375____DOLLAR__1237 ) == ( 8'd2 )  ;
assign n390____DOLLAR__1244 =  ( n375____DOLLAR__1237 ) == ( 8'd1 )  ;
assign n391____DOLLAR__1246 =  ( n390____DOLLAR__1244 ) ? ( 32'd498536548 ) : ( 32'd0 ) ;
assign n392____DOLLAR__1253 =  ( n389____DOLLAR__1251 ) ? ( 32'd997073096 ) : ( n391____DOLLAR__1246 ) ;
assign n393____DOLLAR__1260 =  ( n388____DOLLAR__1258 ) ? ( 32'd651767980 ) : ( n392____DOLLAR__1253 ) ;
assign n394____DOLLAR__1267 =  ( n387____DOLLAR__1265 ) ? ( 32'd1994146192 ) : ( n393____DOLLAR__1260 ) ;
assign n395____DOLLAR__1274 =  ( n386____DOLLAR__1272 ) ? ( 32'd1802195444 ) : ( n394____DOLLAR__1267 ) ;
assign n396____DOLLAR__1281 =  ( n385____DOLLAR__1279 ) ? ( 32'd1303535960 ) : ( n395____DOLLAR__1274 ) ;
assign n397____DOLLAR__1288 =  ( n384____DOLLAR__1286 ) ? ( 32'd1342533948 ) : ( n396____DOLLAR__1281 ) ;
assign n398____DOLLAR__1295 =  ( n383____DOLLAR__1293 ) ? ( 32'd-306674912 ) : ( n397____DOLLAR__1288 ) ;
assign n399____DOLLAR__1302 =  ( n382____DOLLAR__1300 ) ? ( 32'd-267414716 ) : ( n398____DOLLAR__1295 ) ;
assign n400____DOLLAR__1309 =  ( n381____DOLLAR__1307 ) ? ( 32'd-690576408 ) : ( n399____DOLLAR__1302 ) ;
assign n401____DOLLAR__1316 =  ( n380____DOLLAR__1314 ) ? ( 32'd-882789492 ) : ( n400____DOLLAR__1309 ) ;
assign n402____DOLLAR__1323 =  ( n379____DOLLAR__1321 ) ? ( 32'd-1687895376 ) : ( n401____DOLLAR__1316 ) ;
assign n403____DOLLAR__1330 =  ( n378____DOLLAR__1328 ) ? ( 32'd-2032938284 ) : ( n402____DOLLAR__1323 ) ;
assign n404____DOLLAR__1337 =  ( n377____DOLLAR__1335 ) ? ( 32'd-1609899400 ) : ( n403____DOLLAR__1330 ) ;
assign n405____DOLLAR__1344 =  ( n376____DOLLAR__1342 ) ? ( 32'd-1111625188 ) : ( n404____DOLLAR__1337 ) ;
assign n406____DOLLAR__1231 =  ( $signed( n371____DOLLAR__1226 ) >>> ( 32'd4 ))  ;
assign n407____DOLLAR__1345 =  ( n405____DOLLAR__1344 ) ^ ( n406____DOLLAR__1231 )  ;
assign n408____DOLLAR__1354 = n407____DOLLAR__1345[7:0] ;
assign n409____DOLLAR__1353 =  ( $signed( n373____DOLLAR__1227 ) >>> ( 8'd4 ))  ;
assign n410____DOLLAR__1356 =  ( n408____DOLLAR__1354 ) ^ ( n409____DOLLAR__1353 )  ;
assign n411____DOLLAR__1357 =  ( n410____DOLLAR__1356 ) & ( 8'd15 )  ;
assign n412____DOLLAR__1462 =  ( n411____DOLLAR__1357 ) == ( 8'd15 )  ;
assign n413____DOLLAR__1455 =  ( n411____DOLLAR__1357 ) == ( 8'd14 )  ;
assign n414____DOLLAR__1448 =  ( n411____DOLLAR__1357 ) == ( 8'd13 )  ;
assign n415____DOLLAR__1441 =  ( n411____DOLLAR__1357 ) == ( 8'd12 )  ;
assign n416____DOLLAR__1434 =  ( n411____DOLLAR__1357 ) == ( 8'd11 )  ;
assign n417____DOLLAR__1427 =  ( n411____DOLLAR__1357 ) == ( 8'd10 )  ;
assign n418____DOLLAR__1420 =  ( n411____DOLLAR__1357 ) == ( 8'd9 )  ;
assign n419____DOLLAR__1413 =  ( n411____DOLLAR__1357 ) == ( 8'd8 )  ;
assign n420____DOLLAR__1406 =  ( n411____DOLLAR__1357 ) == ( 8'd7 )  ;
assign n421____DOLLAR__1399 =  ( n411____DOLLAR__1357 ) == ( 8'd6 )  ;
assign n422____DOLLAR__1392 =  ( n411____DOLLAR__1357 ) == ( 8'd5 )  ;
assign n423____DOLLAR__1385 =  ( n411____DOLLAR__1357 ) == ( 8'd4 )  ;
assign n424____DOLLAR__1378 =  ( n411____DOLLAR__1357 ) == ( 8'd3 )  ;
assign n425____DOLLAR__1371 =  ( n411____DOLLAR__1357 ) == ( 8'd2 )  ;
assign n426____DOLLAR__1364 =  ( n411____DOLLAR__1357 ) == ( 8'd1 )  ;
assign n427____DOLLAR__1366 =  ( n426____DOLLAR__1364 ) ? ( 32'd498536548 ) : ( 32'd0 ) ;
assign n428____DOLLAR__1373 =  ( n425____DOLLAR__1371 ) ? ( 32'd997073096 ) : ( n427____DOLLAR__1366 ) ;
assign n429____DOLLAR__1380 =  ( n424____DOLLAR__1378 ) ? ( 32'd651767980 ) : ( n428____DOLLAR__1373 ) ;
assign n430____DOLLAR__1387 =  ( n423____DOLLAR__1385 ) ? ( 32'd1994146192 ) : ( n429____DOLLAR__1380 ) ;
assign n431____DOLLAR__1394 =  ( n422____DOLLAR__1392 ) ? ( 32'd1802195444 ) : ( n430____DOLLAR__1387 ) ;
assign n432____DOLLAR__1401 =  ( n421____DOLLAR__1399 ) ? ( 32'd1303535960 ) : ( n431____DOLLAR__1394 ) ;
assign n433____DOLLAR__1408 =  ( n420____DOLLAR__1406 ) ? ( 32'd1342533948 ) : ( n432____DOLLAR__1401 ) ;
assign n434____DOLLAR__1415 =  ( n419____DOLLAR__1413 ) ? ( 32'd-306674912 ) : ( n433____DOLLAR__1408 ) ;
assign n435____DOLLAR__1422 =  ( n418____DOLLAR__1420 ) ? ( 32'd-267414716 ) : ( n434____DOLLAR__1415 ) ;
assign n436____DOLLAR__1429 =  ( n417____DOLLAR__1427 ) ? ( 32'd-690576408 ) : ( n435____DOLLAR__1422 ) ;
assign n437____DOLLAR__1436 =  ( n416____DOLLAR__1434 ) ? ( 32'd-882789492 ) : ( n436____DOLLAR__1429 ) ;
assign n438____DOLLAR__1443 =  ( n415____DOLLAR__1441 ) ? ( 32'd-1687895376 ) : ( n437____DOLLAR__1436 ) ;
assign n439____DOLLAR__1450 =  ( n414____DOLLAR__1448 ) ? ( 32'd-2032938284 ) : ( n438____DOLLAR__1443 ) ;
assign n440____DOLLAR__1457 =  ( n413____DOLLAR__1455 ) ? ( 32'd-1609899400 ) : ( n439____DOLLAR__1450 ) ;
assign n441____DOLLAR__1464 =  ( n412____DOLLAR__1462 ) ? ( 32'd-1111625188 ) : ( n440____DOLLAR__1457 ) ;
assign n442____DOLLAR__1348 =  ( $signed( n407____DOLLAR__1345 ) >>> ( 32'd4 ))  ;
assign n443____DOLLAR__1465 =  ( n441____DOLLAR__1464 ) ^ ( n442____DOLLAR__1348 )  ;
assign n444____DOLLAR__1473 = n443____DOLLAR__1465[7:0] ;
assign n445____DOLLAR__1466 = CRC_DAT_IN[31:24] ;
assign n446____DOLLAR__1475 =  ( n444____DOLLAR__1473 ) ^ ( n445____DOLLAR__1466 )  ;
assign n447____DOLLAR__1476 =  ( n446____DOLLAR__1475 ) & ( 8'd15 )  ;
assign n448____DOLLAR__1581 =  ( n447____DOLLAR__1476 ) == ( 8'd15 )  ;
assign n449____DOLLAR__1574 =  ( n447____DOLLAR__1476 ) == ( 8'd14 )  ;
assign n450____DOLLAR__1567 =  ( n447____DOLLAR__1476 ) == ( 8'd13 )  ;
assign n451____DOLLAR__1560 =  ( n447____DOLLAR__1476 ) == ( 8'd12 )  ;
assign n452____DOLLAR__1553 =  ( n447____DOLLAR__1476 ) == ( 8'd11 )  ;
assign n453____DOLLAR__1546 =  ( n447____DOLLAR__1476 ) == ( 8'd10 )  ;
assign n454____DOLLAR__1539 =  ( n447____DOLLAR__1476 ) == ( 8'd9 )  ;
assign n455____DOLLAR__1532 =  ( n447____DOLLAR__1476 ) == ( 8'd8 )  ;
assign n456____DOLLAR__1525 =  ( n447____DOLLAR__1476 ) == ( 8'd7 )  ;
assign n457____DOLLAR__1518 =  ( n447____DOLLAR__1476 ) == ( 8'd6 )  ;
assign n458____DOLLAR__1511 =  ( n447____DOLLAR__1476 ) == ( 8'd5 )  ;
assign n459____DOLLAR__1504 =  ( n447____DOLLAR__1476 ) == ( 8'd4 )  ;
assign n460____DOLLAR__1497 =  ( n447____DOLLAR__1476 ) == ( 8'd3 )  ;
assign n461____DOLLAR__1490 =  ( n447____DOLLAR__1476 ) == ( 8'd2 )  ;
assign n462____DOLLAR__1483 =  ( n447____DOLLAR__1476 ) == ( 8'd1 )  ;
assign n463____DOLLAR__1485 =  ( n462____DOLLAR__1483 ) ? ( 32'd498536548 ) : ( 32'd0 ) ;
assign n464____DOLLAR__1492 =  ( n461____DOLLAR__1490 ) ? ( 32'd997073096 ) : ( n463____DOLLAR__1485 ) ;
assign n465____DOLLAR__1499 =  ( n460____DOLLAR__1497 ) ? ( 32'd651767980 ) : ( n464____DOLLAR__1492 ) ;
assign n466____DOLLAR__1506 =  ( n459____DOLLAR__1504 ) ? ( 32'd1994146192 ) : ( n465____DOLLAR__1499 ) ;
assign n467____DOLLAR__1513 =  ( n458____DOLLAR__1511 ) ? ( 32'd1802195444 ) : ( n466____DOLLAR__1506 ) ;
assign n468____DOLLAR__1520 =  ( n457____DOLLAR__1518 ) ? ( 32'd1303535960 ) : ( n467____DOLLAR__1513 ) ;
assign n469____DOLLAR__1527 =  ( n456____DOLLAR__1525 ) ? ( 32'd1342533948 ) : ( n468____DOLLAR__1520 ) ;
assign n470____DOLLAR__1534 =  ( n455____DOLLAR__1532 ) ? ( 32'd-306674912 ) : ( n469____DOLLAR__1527 ) ;
assign n471____DOLLAR__1541 =  ( n454____DOLLAR__1539 ) ? ( 32'd-267414716 ) : ( n470____DOLLAR__1534 ) ;
assign n472____DOLLAR__1548 =  ( n453____DOLLAR__1546 ) ? ( 32'd-690576408 ) : ( n471____DOLLAR__1541 ) ;
assign n473____DOLLAR__1555 =  ( n452____DOLLAR__1553 ) ? ( 32'd-882789492 ) : ( n472____DOLLAR__1548 ) ;
assign n474____DOLLAR__1562 =  ( n451____DOLLAR__1560 ) ? ( 32'd-1687895376 ) : ( n473____DOLLAR__1555 ) ;
assign n475____DOLLAR__1569 =  ( n450____DOLLAR__1567 ) ? ( 32'd-2032938284 ) : ( n474____DOLLAR__1562 ) ;
assign n476____DOLLAR__1576 =  ( n449____DOLLAR__1574 ) ? ( 32'd-1609899400 ) : ( n475____DOLLAR__1569 ) ;
assign n477____DOLLAR__1583 =  ( n448____DOLLAR__1581 ) ? ( 32'd-1111625188 ) : ( n476____DOLLAR__1576 ) ;
assign n478____DOLLAR__1470 =  ( $signed( n443____DOLLAR__1465 ) >>> ( 32'd4 ))  ;
assign n479____DOLLAR__1584 =  ( n477____DOLLAR__1583 ) ^ ( n478____DOLLAR__1470 )  ;
assign n480____DOLLAR__1593 = n479____DOLLAR__1584[7:0] ;
assign n481____DOLLAR__1592 =  ( $signed( n445____DOLLAR__1466 ) >>> ( 8'd4 ))  ;
assign n482____DOLLAR__1595 =  ( n480____DOLLAR__1593 ) ^ ( n481____DOLLAR__1592 )  ;
assign n483____DOLLAR__1596 =  ( n482____DOLLAR__1595 ) & ( 8'd15 )  ;
assign n484____DOLLAR__1701 =  ( n483____DOLLAR__1596 ) == ( 8'd15 )  ;
assign n485____DOLLAR__1694 =  ( n483____DOLLAR__1596 ) == ( 8'd14 )  ;
assign n486____DOLLAR__1687 =  ( n483____DOLLAR__1596 ) == ( 8'd13 )  ;
assign n487____DOLLAR__1680 =  ( n483____DOLLAR__1596 ) == ( 8'd12 )  ;
assign n488____DOLLAR__1673 =  ( n483____DOLLAR__1596 ) == ( 8'd11 )  ;
assign n489____DOLLAR__1666 =  ( n483____DOLLAR__1596 ) == ( 8'd10 )  ;
assign n490____DOLLAR__1659 =  ( n483____DOLLAR__1596 ) == ( 8'd9 )  ;
assign n491____DOLLAR__1652 =  ( n483____DOLLAR__1596 ) == ( 8'd8 )  ;
assign n492____DOLLAR__1645 =  ( n483____DOLLAR__1596 ) == ( 8'd7 )  ;
assign n493____DOLLAR__1638 =  ( n483____DOLLAR__1596 ) == ( 8'd6 )  ;
assign n494____DOLLAR__1631 =  ( n483____DOLLAR__1596 ) == ( 8'd5 )  ;
assign n495____DOLLAR__1624 =  ( n483____DOLLAR__1596 ) == ( 8'd4 )  ;
assign n496____DOLLAR__1617 =  ( n483____DOLLAR__1596 ) == ( 8'd3 )  ;
assign n497____DOLLAR__1610 =  ( n483____DOLLAR__1596 ) == ( 8'd2 )  ;
assign n498____DOLLAR__1603 =  ( n483____DOLLAR__1596 ) == ( 8'd1 )  ;
assign n499____DOLLAR__1605 =  ( n498____DOLLAR__1603 ) ? ( 32'd498536548 ) : ( 32'd0 ) ;
assign n500____DOLLAR__1612 =  ( n497____DOLLAR__1610 ) ? ( 32'd997073096 ) : ( n499____DOLLAR__1605 ) ;
assign n501____DOLLAR__1619 =  ( n496____DOLLAR__1617 ) ? ( 32'd651767980 ) : ( n500____DOLLAR__1612 ) ;
assign n502____DOLLAR__1626 =  ( n495____DOLLAR__1624 ) ? ( 32'd1994146192 ) : ( n501____DOLLAR__1619 ) ;
assign n503____DOLLAR__1633 =  ( n494____DOLLAR__1631 ) ? ( 32'd1802195444 ) : ( n502____DOLLAR__1626 ) ;
assign n504____DOLLAR__1640 =  ( n493____DOLLAR__1638 ) ? ( 32'd1303535960 ) : ( n503____DOLLAR__1633 ) ;
assign n505____DOLLAR__1647 =  ( n492____DOLLAR__1645 ) ? ( 32'd1342533948 ) : ( n504____DOLLAR__1640 ) ;
assign n506____DOLLAR__1654 =  ( n491____DOLLAR__1652 ) ? ( 32'd-306674912 ) : ( n505____DOLLAR__1647 ) ;
assign n507____DOLLAR__1661 =  ( n490____DOLLAR__1659 ) ? ( 32'd-267414716 ) : ( n506____DOLLAR__1654 ) ;
assign n508____DOLLAR__1668 =  ( n489____DOLLAR__1666 ) ? ( 32'd-690576408 ) : ( n507____DOLLAR__1661 ) ;
assign n509____DOLLAR__1675 =  ( n488____DOLLAR__1673 ) ? ( 32'd-882789492 ) : ( n508____DOLLAR__1668 ) ;
assign n510____DOLLAR__1682 =  ( n487____DOLLAR__1680 ) ? ( 32'd-1687895376 ) : ( n509____DOLLAR__1675 ) ;
assign n511____DOLLAR__1689 =  ( n486____DOLLAR__1687 ) ? ( 32'd-2032938284 ) : ( n510____DOLLAR__1682 ) ;
assign n512____DOLLAR__1696 =  ( n485____DOLLAR__1694 ) ? ( 32'd-1609899400 ) : ( n511____DOLLAR__1689 ) ;
assign n513____DOLLAR__1703 =  ( n484____DOLLAR__1701 ) ? ( 32'd-1111625188 ) : ( n512____DOLLAR__1696 ) ;
assign n514____DOLLAR__1587 =  ( $signed( n479____DOLLAR__1584 ) >>> ( 32'd4 ))  ;
assign n515____DOLLAR__1704 =  ( n513____DOLLAR__1703 ) ^ ( n514____DOLLAR__1587 )  ;
assign n516____DOLLAR__1712 = n515____DOLLAR__1704[7:0] ;
assign n517____DOLLAR__1705 = CRC_DAT_IN[39:32] ;
assign n518____DOLLAR__1714 =  ( n516____DOLLAR__1712 ) ^ ( n517____DOLLAR__1705 )  ;
assign n519____DOLLAR__1715 =  ( n518____DOLLAR__1714 ) & ( 8'd15 )  ;
assign n520____DOLLAR__1820 =  ( n519____DOLLAR__1715 ) == ( 8'd15 )  ;
assign n521____DOLLAR__1813 =  ( n519____DOLLAR__1715 ) == ( 8'd14 )  ;
assign n522____DOLLAR__1806 =  ( n519____DOLLAR__1715 ) == ( 8'd13 )  ;
assign n523____DOLLAR__1799 =  ( n519____DOLLAR__1715 ) == ( 8'd12 )  ;
assign n524____DOLLAR__1792 =  ( n519____DOLLAR__1715 ) == ( 8'd11 )  ;
assign n525____DOLLAR__1785 =  ( n519____DOLLAR__1715 ) == ( 8'd10 )  ;
assign n526____DOLLAR__1778 =  ( n519____DOLLAR__1715 ) == ( 8'd9 )  ;
assign n527____DOLLAR__1771 =  ( n519____DOLLAR__1715 ) == ( 8'd8 )  ;
assign n528____DOLLAR__1764 =  ( n519____DOLLAR__1715 ) == ( 8'd7 )  ;
assign n529____DOLLAR__1757 =  ( n519____DOLLAR__1715 ) == ( 8'd6 )  ;
assign n530____DOLLAR__1750 =  ( n519____DOLLAR__1715 ) == ( 8'd5 )  ;
assign n531____DOLLAR__1743 =  ( n519____DOLLAR__1715 ) == ( 8'd4 )  ;
assign n532____DOLLAR__1736 =  ( n519____DOLLAR__1715 ) == ( 8'd3 )  ;
assign n533____DOLLAR__1729 =  ( n519____DOLLAR__1715 ) == ( 8'd2 )  ;
assign n534____DOLLAR__1722 =  ( n519____DOLLAR__1715 ) == ( 8'd1 )  ;
assign n535____DOLLAR__1724 =  ( n534____DOLLAR__1722 ) ? ( 32'd498536548 ) : ( 32'd0 ) ;
assign n536____DOLLAR__1731 =  ( n533____DOLLAR__1729 ) ? ( 32'd997073096 ) : ( n535____DOLLAR__1724 ) ;
assign n537____DOLLAR__1738 =  ( n532____DOLLAR__1736 ) ? ( 32'd651767980 ) : ( n536____DOLLAR__1731 ) ;
assign n538____DOLLAR__1745 =  ( n531____DOLLAR__1743 ) ? ( 32'd1994146192 ) : ( n537____DOLLAR__1738 ) ;
assign n539____DOLLAR__1752 =  ( n530____DOLLAR__1750 ) ? ( 32'd1802195444 ) : ( n538____DOLLAR__1745 ) ;
assign n540____DOLLAR__1759 =  ( n529____DOLLAR__1757 ) ? ( 32'd1303535960 ) : ( n539____DOLLAR__1752 ) ;
assign n541____DOLLAR__1766 =  ( n528____DOLLAR__1764 ) ? ( 32'd1342533948 ) : ( n540____DOLLAR__1759 ) ;
assign n542____DOLLAR__1773 =  ( n527____DOLLAR__1771 ) ? ( 32'd-306674912 ) : ( n541____DOLLAR__1766 ) ;
assign n543____DOLLAR__1780 =  ( n526____DOLLAR__1778 ) ? ( 32'd-267414716 ) : ( n542____DOLLAR__1773 ) ;
assign n544____DOLLAR__1787 =  ( n525____DOLLAR__1785 ) ? ( 32'd-690576408 ) : ( n543____DOLLAR__1780 ) ;
assign n545____DOLLAR__1794 =  ( n524____DOLLAR__1792 ) ? ( 32'd-882789492 ) : ( n544____DOLLAR__1787 ) ;
assign n546____DOLLAR__1801 =  ( n523____DOLLAR__1799 ) ? ( 32'd-1687895376 ) : ( n545____DOLLAR__1794 ) ;
assign n547____DOLLAR__1808 =  ( n522____DOLLAR__1806 ) ? ( 32'd-2032938284 ) : ( n546____DOLLAR__1801 ) ;
assign n548____DOLLAR__1815 =  ( n521____DOLLAR__1813 ) ? ( 32'd-1609899400 ) : ( n547____DOLLAR__1808 ) ;
assign n549____DOLLAR__1822 =  ( n520____DOLLAR__1820 ) ? ( 32'd-1111625188 ) : ( n548____DOLLAR__1815 ) ;
assign n550____DOLLAR__1709 =  ( $signed( n515____DOLLAR__1704 ) >>> ( 32'd4 ))  ;
assign n551____DOLLAR__1823 =  ( n549____DOLLAR__1822 ) ^ ( n550____DOLLAR__1709 )  ;
assign n552____DOLLAR__1832 = n551____DOLLAR__1823[7:0] ;
assign n553____DOLLAR__1831 =  ( $signed( n517____DOLLAR__1705 ) >>> ( 8'd4 ))  ;
assign n554____DOLLAR__1834 =  ( n552____DOLLAR__1832 ) ^ ( n553____DOLLAR__1831 )  ;
assign n555____DOLLAR__1835 =  ( n554____DOLLAR__1834 ) & ( 8'd15 )  ;
assign n556____DOLLAR__1940 =  ( n555____DOLLAR__1835 ) == ( 8'd15 )  ;
assign n557____DOLLAR__1933 =  ( n555____DOLLAR__1835 ) == ( 8'd14 )  ;
assign n558____DOLLAR__1926 =  ( n555____DOLLAR__1835 ) == ( 8'd13 )  ;
assign n559____DOLLAR__1919 =  ( n555____DOLLAR__1835 ) == ( 8'd12 )  ;
assign n560____DOLLAR__1912 =  ( n555____DOLLAR__1835 ) == ( 8'd11 )  ;
assign n561____DOLLAR__1905 =  ( n555____DOLLAR__1835 ) == ( 8'd10 )  ;
assign n562____DOLLAR__1898 =  ( n555____DOLLAR__1835 ) == ( 8'd9 )  ;
assign n563____DOLLAR__1891 =  ( n555____DOLLAR__1835 ) == ( 8'd8 )  ;
assign n564____DOLLAR__1884 =  ( n555____DOLLAR__1835 ) == ( 8'd7 )  ;
assign n565____DOLLAR__1877 =  ( n555____DOLLAR__1835 ) == ( 8'd6 )  ;
assign n566____DOLLAR__1870 =  ( n555____DOLLAR__1835 ) == ( 8'd5 )  ;
assign n567____DOLLAR__1863 =  ( n555____DOLLAR__1835 ) == ( 8'd4 )  ;
assign n568____DOLLAR__1856 =  ( n555____DOLLAR__1835 ) == ( 8'd3 )  ;
assign n569____DOLLAR__1849 =  ( n555____DOLLAR__1835 ) == ( 8'd2 )  ;
assign n570____DOLLAR__1842 =  ( n555____DOLLAR__1835 ) == ( 8'd1 )  ;
assign n571____DOLLAR__1844 =  ( n570____DOLLAR__1842 ) ? ( 32'd498536548 ) : ( 32'd0 ) ;
assign n572____DOLLAR__1851 =  ( n569____DOLLAR__1849 ) ? ( 32'd997073096 ) : ( n571____DOLLAR__1844 ) ;
assign n573____DOLLAR__1858 =  ( n568____DOLLAR__1856 ) ? ( 32'd651767980 ) : ( n572____DOLLAR__1851 ) ;
assign n574____DOLLAR__1865 =  ( n567____DOLLAR__1863 ) ? ( 32'd1994146192 ) : ( n573____DOLLAR__1858 ) ;
assign n575____DOLLAR__1872 =  ( n566____DOLLAR__1870 ) ? ( 32'd1802195444 ) : ( n574____DOLLAR__1865 ) ;
assign n576____DOLLAR__1879 =  ( n565____DOLLAR__1877 ) ? ( 32'd1303535960 ) : ( n575____DOLLAR__1872 ) ;
assign n577____DOLLAR__1886 =  ( n564____DOLLAR__1884 ) ? ( 32'd1342533948 ) : ( n576____DOLLAR__1879 ) ;
assign n578____DOLLAR__1893 =  ( n563____DOLLAR__1891 ) ? ( 32'd-306674912 ) : ( n577____DOLLAR__1886 ) ;
assign n579____DOLLAR__1900 =  ( n562____DOLLAR__1898 ) ? ( 32'd-267414716 ) : ( n578____DOLLAR__1893 ) ;
assign n580____DOLLAR__1907 =  ( n561____DOLLAR__1905 ) ? ( 32'd-690576408 ) : ( n579____DOLLAR__1900 ) ;
assign n581____DOLLAR__1914 =  ( n560____DOLLAR__1912 ) ? ( 32'd-882789492 ) : ( n580____DOLLAR__1907 ) ;
assign n582____DOLLAR__1921 =  ( n559____DOLLAR__1919 ) ? ( 32'd-1687895376 ) : ( n581____DOLLAR__1914 ) ;
assign n583____DOLLAR__1928 =  ( n558____DOLLAR__1926 ) ? ( 32'd-2032938284 ) : ( n582____DOLLAR__1921 ) ;
assign n584____DOLLAR__1935 =  ( n557____DOLLAR__1933 ) ? ( 32'd-1609899400 ) : ( n583____DOLLAR__1928 ) ;
assign n585____DOLLAR__1942 =  ( n556____DOLLAR__1940 ) ? ( 32'd-1111625188 ) : ( n584____DOLLAR__1935 ) ;
assign n586____DOLLAR__1826 =  ( $signed( n551____DOLLAR__1823 ) >>> ( 32'd4 ))  ;
assign n587____DOLLAR__1943 =  ( n585____DOLLAR__1942 ) ^ ( n586____DOLLAR__1826 )  ;
assign n588____DOLLAR__1951 = n587____DOLLAR__1943[7:0] ;
assign n589____DOLLAR__1944 = CRC_DAT_IN[47:40] ;
assign n590____DOLLAR__1953 =  ( n588____DOLLAR__1951 ) ^ ( n589____DOLLAR__1944 )  ;
assign n591____DOLLAR__1954 =  ( n590____DOLLAR__1953 ) & ( 8'd15 )  ;
assign n592____DOLLAR__2059 =  ( n591____DOLLAR__1954 ) == ( 8'd15 )  ;
assign n593____DOLLAR__2052 =  ( n591____DOLLAR__1954 ) == ( 8'd14 )  ;
assign n594____DOLLAR__2045 =  ( n591____DOLLAR__1954 ) == ( 8'd13 )  ;
assign n595____DOLLAR__2038 =  ( n591____DOLLAR__1954 ) == ( 8'd12 )  ;
assign n596____DOLLAR__2031 =  ( n591____DOLLAR__1954 ) == ( 8'd11 )  ;
assign n597____DOLLAR__2024 =  ( n591____DOLLAR__1954 ) == ( 8'd10 )  ;
assign n598____DOLLAR__2017 =  ( n591____DOLLAR__1954 ) == ( 8'd9 )  ;
assign n599____DOLLAR__2010 =  ( n591____DOLLAR__1954 ) == ( 8'd8 )  ;
assign n600____DOLLAR__2003 =  ( n591____DOLLAR__1954 ) == ( 8'd7 )  ;
assign n601____DOLLAR__1996 =  ( n591____DOLLAR__1954 ) == ( 8'd6 )  ;
assign n602____DOLLAR__1989 =  ( n591____DOLLAR__1954 ) == ( 8'd5 )  ;
assign n603____DOLLAR__1982 =  ( n591____DOLLAR__1954 ) == ( 8'd4 )  ;
assign n604____DOLLAR__1975 =  ( n591____DOLLAR__1954 ) == ( 8'd3 )  ;
assign n605____DOLLAR__1968 =  ( n591____DOLLAR__1954 ) == ( 8'd2 )  ;
assign n606____DOLLAR__1961 =  ( n591____DOLLAR__1954 ) == ( 8'd1 )  ;
assign n607____DOLLAR__1963 =  ( n606____DOLLAR__1961 ) ? ( 32'd498536548 ) : ( 32'd0 ) ;
assign n608____DOLLAR__1970 =  ( n605____DOLLAR__1968 ) ? ( 32'd997073096 ) : ( n607____DOLLAR__1963 ) ;
assign n609____DOLLAR__1977 =  ( n604____DOLLAR__1975 ) ? ( 32'd651767980 ) : ( n608____DOLLAR__1970 ) ;
assign n610____DOLLAR__1984 =  ( n603____DOLLAR__1982 ) ? ( 32'd1994146192 ) : ( n609____DOLLAR__1977 ) ;
assign n611____DOLLAR__1991 =  ( n602____DOLLAR__1989 ) ? ( 32'd1802195444 ) : ( n610____DOLLAR__1984 ) ;
assign n612____DOLLAR__1998 =  ( n601____DOLLAR__1996 ) ? ( 32'd1303535960 ) : ( n611____DOLLAR__1991 ) ;
assign n613____DOLLAR__2005 =  ( n600____DOLLAR__2003 ) ? ( 32'd1342533948 ) : ( n612____DOLLAR__1998 ) ;
assign n614____DOLLAR__2012 =  ( n599____DOLLAR__2010 ) ? ( 32'd-306674912 ) : ( n613____DOLLAR__2005 ) ;
assign n615____DOLLAR__2019 =  ( n598____DOLLAR__2017 ) ? ( 32'd-267414716 ) : ( n614____DOLLAR__2012 ) ;
assign n616____DOLLAR__2026 =  ( n597____DOLLAR__2024 ) ? ( 32'd-690576408 ) : ( n615____DOLLAR__2019 ) ;
assign n617____DOLLAR__2033 =  ( n596____DOLLAR__2031 ) ? ( 32'd-882789492 ) : ( n616____DOLLAR__2026 ) ;
assign n618____DOLLAR__2040 =  ( n595____DOLLAR__2038 ) ? ( 32'd-1687895376 ) : ( n617____DOLLAR__2033 ) ;
assign n619____DOLLAR__2047 =  ( n594____DOLLAR__2045 ) ? ( 32'd-2032938284 ) : ( n618____DOLLAR__2040 ) ;
assign n620____DOLLAR__2054 =  ( n593____DOLLAR__2052 ) ? ( 32'd-1609899400 ) : ( n619____DOLLAR__2047 ) ;
assign n621____DOLLAR__2061 =  ( n592____DOLLAR__2059 ) ? ( 32'd-1111625188 ) : ( n620____DOLLAR__2054 ) ;
assign n622____DOLLAR__1948 =  ( $signed( n587____DOLLAR__1943 ) >>> ( 32'd4 ))  ;
assign n623____DOLLAR__2062 =  ( n621____DOLLAR__2061 ) ^ ( n622____DOLLAR__1948 )  ;
assign n624____DOLLAR__2071 = n623____DOLLAR__2062[7:0] ;
assign n625____DOLLAR__2070 =  ( $signed( n589____DOLLAR__1944 ) >>> ( 8'd4 ))  ;
assign n626____DOLLAR__2073 =  ( n624____DOLLAR__2071 ) ^ ( n625____DOLLAR__2070 )  ;
assign n627____DOLLAR__2074 =  ( n626____DOLLAR__2073 ) & ( 8'd15 )  ;
assign n628____DOLLAR__2179 =  ( n627____DOLLAR__2074 ) == ( 8'd15 )  ;
assign n629____DOLLAR__2172 =  ( n627____DOLLAR__2074 ) == ( 8'd14 )  ;
assign n630____DOLLAR__2165 =  ( n627____DOLLAR__2074 ) == ( 8'd13 )  ;
assign n631____DOLLAR__2158 =  ( n627____DOLLAR__2074 ) == ( 8'd12 )  ;
assign n632____DOLLAR__2151 =  ( n627____DOLLAR__2074 ) == ( 8'd11 )  ;
assign n633____DOLLAR__2144 =  ( n627____DOLLAR__2074 ) == ( 8'd10 )  ;
assign n634____DOLLAR__2137 =  ( n627____DOLLAR__2074 ) == ( 8'd9 )  ;
assign n635____DOLLAR__2130 =  ( n627____DOLLAR__2074 ) == ( 8'd8 )  ;
assign n636____DOLLAR__2123 =  ( n627____DOLLAR__2074 ) == ( 8'd7 )  ;
assign n637____DOLLAR__2116 =  ( n627____DOLLAR__2074 ) == ( 8'd6 )  ;
assign n638____DOLLAR__2109 =  ( n627____DOLLAR__2074 ) == ( 8'd5 )  ;
assign n639____DOLLAR__2102 =  ( n627____DOLLAR__2074 ) == ( 8'd4 )  ;
assign n640____DOLLAR__2095 =  ( n627____DOLLAR__2074 ) == ( 8'd3 )  ;
assign n641____DOLLAR__2088 =  ( n627____DOLLAR__2074 ) == ( 8'd2 )  ;
assign n642____DOLLAR__2081 =  ( n627____DOLLAR__2074 ) == ( 8'd1 )  ;
assign n643____DOLLAR__2083 =  ( n642____DOLLAR__2081 ) ? ( 32'd498536548 ) : ( 32'd0 ) ;
assign n644____DOLLAR__2090 =  ( n641____DOLLAR__2088 ) ? ( 32'd997073096 ) : ( n643____DOLLAR__2083 ) ;
assign n645____DOLLAR__2097 =  ( n640____DOLLAR__2095 ) ? ( 32'd651767980 ) : ( n644____DOLLAR__2090 ) ;
assign n646____DOLLAR__2104 =  ( n639____DOLLAR__2102 ) ? ( 32'd1994146192 ) : ( n645____DOLLAR__2097 ) ;
assign n647____DOLLAR__2111 =  ( n638____DOLLAR__2109 ) ? ( 32'd1802195444 ) : ( n646____DOLLAR__2104 ) ;
assign n648____DOLLAR__2118 =  ( n637____DOLLAR__2116 ) ? ( 32'd1303535960 ) : ( n647____DOLLAR__2111 ) ;
assign n649____DOLLAR__2125 =  ( n636____DOLLAR__2123 ) ? ( 32'd1342533948 ) : ( n648____DOLLAR__2118 ) ;
assign n650____DOLLAR__2132 =  ( n635____DOLLAR__2130 ) ? ( 32'd-306674912 ) : ( n649____DOLLAR__2125 ) ;
assign n651____DOLLAR__2139 =  ( n634____DOLLAR__2137 ) ? ( 32'd-267414716 ) : ( n650____DOLLAR__2132 ) ;
assign n652____DOLLAR__2146 =  ( n633____DOLLAR__2144 ) ? ( 32'd-690576408 ) : ( n651____DOLLAR__2139 ) ;
assign n653____DOLLAR__2153 =  ( n632____DOLLAR__2151 ) ? ( 32'd-882789492 ) : ( n652____DOLLAR__2146 ) ;
assign n654____DOLLAR__2160 =  ( n631____DOLLAR__2158 ) ? ( 32'd-1687895376 ) : ( n653____DOLLAR__2153 ) ;
assign n655____DOLLAR__2167 =  ( n630____DOLLAR__2165 ) ? ( 32'd-2032938284 ) : ( n654____DOLLAR__2160 ) ;
assign n656____DOLLAR__2174 =  ( n629____DOLLAR__2172 ) ? ( 32'd-1609899400 ) : ( n655____DOLLAR__2167 ) ;
assign n657____DOLLAR__2181 =  ( n628____DOLLAR__2179 ) ? ( 32'd-1111625188 ) : ( n656____DOLLAR__2174 ) ;
assign n658____DOLLAR__2065 =  ( $signed( n623____DOLLAR__2062 ) >>> ( 32'd4 ))  ;
assign n659____DOLLAR__2182 =  ( n657____DOLLAR__2181 ) ^ ( n658____DOLLAR__2065 )  ;
assign n660____DOLLAR__2190 = n659____DOLLAR__2182[7:0] ;
assign n661____DOLLAR__2183 = CRC_DAT_IN[55:48] ;
assign n662____DOLLAR__2192 =  ( n660____DOLLAR__2190 ) ^ ( n661____DOLLAR__2183 )  ;
assign n663____DOLLAR__2193 =  ( n662____DOLLAR__2192 ) & ( 8'd15 )  ;
assign n664____DOLLAR__2298 =  ( n663____DOLLAR__2193 ) == ( 8'd15 )  ;
assign n665____DOLLAR__2291 =  ( n663____DOLLAR__2193 ) == ( 8'd14 )  ;
assign n666____DOLLAR__2284 =  ( n663____DOLLAR__2193 ) == ( 8'd13 )  ;
assign n667____DOLLAR__2277 =  ( n663____DOLLAR__2193 ) == ( 8'd12 )  ;
assign n668____DOLLAR__2270 =  ( n663____DOLLAR__2193 ) == ( 8'd11 )  ;
assign n669____DOLLAR__2263 =  ( n663____DOLLAR__2193 ) == ( 8'd10 )  ;
assign n670____DOLLAR__2256 =  ( n663____DOLLAR__2193 ) == ( 8'd9 )  ;
assign n671____DOLLAR__2249 =  ( n663____DOLLAR__2193 ) == ( 8'd8 )  ;
assign n672____DOLLAR__2242 =  ( n663____DOLLAR__2193 ) == ( 8'd7 )  ;
assign n673____DOLLAR__2235 =  ( n663____DOLLAR__2193 ) == ( 8'd6 )  ;
assign n674____DOLLAR__2228 =  ( n663____DOLLAR__2193 ) == ( 8'd5 )  ;
assign n675____DOLLAR__2221 =  ( n663____DOLLAR__2193 ) == ( 8'd4 )  ;
assign n676____DOLLAR__2214 =  ( n663____DOLLAR__2193 ) == ( 8'd3 )  ;
assign n677____DOLLAR__2207 =  ( n663____DOLLAR__2193 ) == ( 8'd2 )  ;
assign n678____DOLLAR__2200 =  ( n663____DOLLAR__2193 ) == ( 8'd1 )  ;
assign n679____DOLLAR__2202 =  ( n678____DOLLAR__2200 ) ? ( 32'd498536548 ) : ( 32'd0 ) ;
assign n680____DOLLAR__2209 =  ( n677____DOLLAR__2207 ) ? ( 32'd997073096 ) : ( n679____DOLLAR__2202 ) ;
assign n681____DOLLAR__2216 =  ( n676____DOLLAR__2214 ) ? ( 32'd651767980 ) : ( n680____DOLLAR__2209 ) ;
assign n682____DOLLAR__2223 =  ( n675____DOLLAR__2221 ) ? ( 32'd1994146192 ) : ( n681____DOLLAR__2216 ) ;
assign n683____DOLLAR__2230 =  ( n674____DOLLAR__2228 ) ? ( 32'd1802195444 ) : ( n682____DOLLAR__2223 ) ;
assign n684____DOLLAR__2237 =  ( n673____DOLLAR__2235 ) ? ( 32'd1303535960 ) : ( n683____DOLLAR__2230 ) ;
assign n685____DOLLAR__2244 =  ( n672____DOLLAR__2242 ) ? ( 32'd1342533948 ) : ( n684____DOLLAR__2237 ) ;
assign n686____DOLLAR__2251 =  ( n671____DOLLAR__2249 ) ? ( 32'd-306674912 ) : ( n685____DOLLAR__2244 ) ;
assign n687____DOLLAR__2258 =  ( n670____DOLLAR__2256 ) ? ( 32'd-267414716 ) : ( n686____DOLLAR__2251 ) ;
assign n688____DOLLAR__2265 =  ( n669____DOLLAR__2263 ) ? ( 32'd-690576408 ) : ( n687____DOLLAR__2258 ) ;
assign n689____DOLLAR__2272 =  ( n668____DOLLAR__2270 ) ? ( 32'd-882789492 ) : ( n688____DOLLAR__2265 ) ;
assign n690____DOLLAR__2279 =  ( n667____DOLLAR__2277 ) ? ( 32'd-1687895376 ) : ( n689____DOLLAR__2272 ) ;
assign n691____DOLLAR__2286 =  ( n666____DOLLAR__2284 ) ? ( 32'd-2032938284 ) : ( n690____DOLLAR__2279 ) ;
assign n692____DOLLAR__2293 =  ( n665____DOLLAR__2291 ) ? ( 32'd-1609899400 ) : ( n691____DOLLAR__2286 ) ;
assign n693____DOLLAR__2300 =  ( n664____DOLLAR__2298 ) ? ( 32'd-1111625188 ) : ( n692____DOLLAR__2293 ) ;
assign n694____DOLLAR__2187 =  ( $signed( n659____DOLLAR__2182 ) >>> ( 32'd4 ))  ;
assign n695____DOLLAR__2301 =  ( n693____DOLLAR__2300 ) ^ ( n694____DOLLAR__2187 )  ;
assign n696____DOLLAR__2310 = n695____DOLLAR__2301[7:0] ;
assign n697____DOLLAR__2309 =  ( $signed( n661____DOLLAR__2183 ) >>> ( 8'd4 ))  ;
assign n698____DOLLAR__2312 =  ( n696____DOLLAR__2310 ) ^ ( n697____DOLLAR__2309 )  ;
assign n699____DOLLAR__2313 =  ( n698____DOLLAR__2312 ) & ( 8'd15 )  ;
assign n700____DOLLAR__2418 =  ( n699____DOLLAR__2313 ) == ( 8'd15 )  ;
assign n701____DOLLAR__2411 =  ( n699____DOLLAR__2313 ) == ( 8'd14 )  ;
assign n702____DOLLAR__2404 =  ( n699____DOLLAR__2313 ) == ( 8'd13 )  ;
assign n703____DOLLAR__2397 =  ( n699____DOLLAR__2313 ) == ( 8'd12 )  ;
assign n704____DOLLAR__2390 =  ( n699____DOLLAR__2313 ) == ( 8'd11 )  ;
assign n705____DOLLAR__2383 =  ( n699____DOLLAR__2313 ) == ( 8'd10 )  ;
assign n706____DOLLAR__2376 =  ( n699____DOLLAR__2313 ) == ( 8'd9 )  ;
assign n707____DOLLAR__2369 =  ( n699____DOLLAR__2313 ) == ( 8'd8 )  ;
assign n708____DOLLAR__2362 =  ( n699____DOLLAR__2313 ) == ( 8'd7 )  ;
assign n709____DOLLAR__2355 =  ( n699____DOLLAR__2313 ) == ( 8'd6 )  ;
assign n710____DOLLAR__2348 =  ( n699____DOLLAR__2313 ) == ( 8'd5 )  ;
assign n711____DOLLAR__2341 =  ( n699____DOLLAR__2313 ) == ( 8'd4 )  ;
assign n712____DOLLAR__2334 =  ( n699____DOLLAR__2313 ) == ( 8'd3 )  ;
assign n713____DOLLAR__2327 =  ( n699____DOLLAR__2313 ) == ( 8'd2 )  ;
assign n714____DOLLAR__2320 =  ( n699____DOLLAR__2313 ) == ( 8'd1 )  ;
assign n715____DOLLAR__2322 =  ( n714____DOLLAR__2320 ) ? ( 32'd498536548 ) : ( 32'd0 ) ;
assign n716____DOLLAR__2329 =  ( n713____DOLLAR__2327 ) ? ( 32'd997073096 ) : ( n715____DOLLAR__2322 ) ;
assign n717____DOLLAR__2336 =  ( n712____DOLLAR__2334 ) ? ( 32'd651767980 ) : ( n716____DOLLAR__2329 ) ;
assign n718____DOLLAR__2343 =  ( n711____DOLLAR__2341 ) ? ( 32'd1994146192 ) : ( n717____DOLLAR__2336 ) ;
assign n719____DOLLAR__2350 =  ( n710____DOLLAR__2348 ) ? ( 32'd1802195444 ) : ( n718____DOLLAR__2343 ) ;
assign n720____DOLLAR__2357 =  ( n709____DOLLAR__2355 ) ? ( 32'd1303535960 ) : ( n719____DOLLAR__2350 ) ;
assign n721____DOLLAR__2364 =  ( n708____DOLLAR__2362 ) ? ( 32'd1342533948 ) : ( n720____DOLLAR__2357 ) ;
assign n722____DOLLAR__2371 =  ( n707____DOLLAR__2369 ) ? ( 32'd-306674912 ) : ( n721____DOLLAR__2364 ) ;
assign n723____DOLLAR__2378 =  ( n706____DOLLAR__2376 ) ? ( 32'd-267414716 ) : ( n722____DOLLAR__2371 ) ;
assign n724____DOLLAR__2385 =  ( n705____DOLLAR__2383 ) ? ( 32'd-690576408 ) : ( n723____DOLLAR__2378 ) ;
assign n725____DOLLAR__2392 =  ( n704____DOLLAR__2390 ) ? ( 32'd-882789492 ) : ( n724____DOLLAR__2385 ) ;
assign n726____DOLLAR__2399 =  ( n703____DOLLAR__2397 ) ? ( 32'd-1687895376 ) : ( n725____DOLLAR__2392 ) ;
assign n727____DOLLAR__2406 =  ( n702____DOLLAR__2404 ) ? ( 32'd-2032938284 ) : ( n726____DOLLAR__2399 ) ;
assign n728____DOLLAR__2413 =  ( n701____DOLLAR__2411 ) ? ( 32'd-1609899400 ) : ( n727____DOLLAR__2406 ) ;
assign n729____DOLLAR__2420 =  ( n700____DOLLAR__2418 ) ? ( 32'd-1111625188 ) : ( n728____DOLLAR__2413 ) ;
assign n730____DOLLAR__2304 =  ( $signed( n695____DOLLAR__2301 ) >>> ( 32'd4 ))  ;
assign n731____DOLLAR__2421 =  ( n729____DOLLAR__2420 ) ^ ( n730____DOLLAR__2304 )  ;
assign n732____DOLLAR__2429 = n731____DOLLAR__2421[7:0] ;
assign n733____DOLLAR__2422 = CRC_DAT_IN[63:56] ;
assign n734____DOLLAR__2431 =  ( n732____DOLLAR__2429 ) ^ ( n733____DOLLAR__2422 )  ;
assign n735____DOLLAR__2432 =  ( n734____DOLLAR__2431 ) & ( 8'd15 )  ;
assign n736____DOLLAR__2537 =  ( n735____DOLLAR__2432 ) == ( 8'd15 )  ;
assign n737____DOLLAR__2530 =  ( n735____DOLLAR__2432 ) == ( 8'd14 )  ;
assign n738____DOLLAR__2523 =  ( n735____DOLLAR__2432 ) == ( 8'd13 )  ;
assign n739____DOLLAR__2516 =  ( n735____DOLLAR__2432 ) == ( 8'd12 )  ;
assign n740____DOLLAR__2509 =  ( n735____DOLLAR__2432 ) == ( 8'd11 )  ;
assign n741____DOLLAR__2502 =  ( n735____DOLLAR__2432 ) == ( 8'd10 )  ;
assign n742____DOLLAR__2495 =  ( n735____DOLLAR__2432 ) == ( 8'd9 )  ;
assign n743____DOLLAR__2488 =  ( n735____DOLLAR__2432 ) == ( 8'd8 )  ;
assign n744____DOLLAR__2481 =  ( n735____DOLLAR__2432 ) == ( 8'd7 )  ;
assign n745____DOLLAR__2474 =  ( n735____DOLLAR__2432 ) == ( 8'd6 )  ;
assign n746____DOLLAR__2467 =  ( n735____DOLLAR__2432 ) == ( 8'd5 )  ;
assign n747____DOLLAR__2460 =  ( n735____DOLLAR__2432 ) == ( 8'd4 )  ;
assign n748____DOLLAR__2453 =  ( n735____DOLLAR__2432 ) == ( 8'd3 )  ;
assign n749____DOLLAR__2446 =  ( n735____DOLLAR__2432 ) == ( 8'd2 )  ;
assign n750____DOLLAR__2439 =  ( n735____DOLLAR__2432 ) == ( 8'd1 )  ;
assign n751____DOLLAR__2441 =  ( n750____DOLLAR__2439 ) ? ( 32'd498536548 ) : ( 32'd0 ) ;
assign n752____DOLLAR__2448 =  ( n749____DOLLAR__2446 ) ? ( 32'd997073096 ) : ( n751____DOLLAR__2441 ) ;
assign n753____DOLLAR__2455 =  ( n748____DOLLAR__2453 ) ? ( 32'd651767980 ) : ( n752____DOLLAR__2448 ) ;
assign n754____DOLLAR__2462 =  ( n747____DOLLAR__2460 ) ? ( 32'd1994146192 ) : ( n753____DOLLAR__2455 ) ;
assign n755____DOLLAR__2469 =  ( n746____DOLLAR__2467 ) ? ( 32'd1802195444 ) : ( n754____DOLLAR__2462 ) ;
assign n756____DOLLAR__2476 =  ( n745____DOLLAR__2474 ) ? ( 32'd1303535960 ) : ( n755____DOLLAR__2469 ) ;
assign n757____DOLLAR__2483 =  ( n744____DOLLAR__2481 ) ? ( 32'd1342533948 ) : ( n756____DOLLAR__2476 ) ;
assign n758____DOLLAR__2490 =  ( n743____DOLLAR__2488 ) ? ( 32'd-306674912 ) : ( n757____DOLLAR__2483 ) ;
assign n759____DOLLAR__2497 =  ( n742____DOLLAR__2495 ) ? ( 32'd-267414716 ) : ( n758____DOLLAR__2490 ) ;
assign n760____DOLLAR__2504 =  ( n741____DOLLAR__2502 ) ? ( 32'd-690576408 ) : ( n759____DOLLAR__2497 ) ;
assign n761____DOLLAR__2511 =  ( n740____DOLLAR__2509 ) ? ( 32'd-882789492 ) : ( n760____DOLLAR__2504 ) ;
assign n762____DOLLAR__2518 =  ( n739____DOLLAR__2516 ) ? ( 32'd-1687895376 ) : ( n761____DOLLAR__2511 ) ;
assign n763____DOLLAR__2525 =  ( n738____DOLLAR__2523 ) ? ( 32'd-2032938284 ) : ( n762____DOLLAR__2518 ) ;
assign n764____DOLLAR__2532 =  ( n737____DOLLAR__2530 ) ? ( 32'd-1609899400 ) : ( n763____DOLLAR__2525 ) ;
assign n765____DOLLAR__2539 =  ( n736____DOLLAR__2537 ) ? ( 32'd-1111625188 ) : ( n764____DOLLAR__2532 ) ;
assign n766____DOLLAR__2426 =  ( $signed( n731____DOLLAR__2421 ) >>> ( 32'd4 ))  ;
assign n767____DOLLAR__2540 =  ( n765____DOLLAR__2539 ) ^ ( n766____DOLLAR__2426 )  ;
assign n768____DOLLAR__2549 = n767____DOLLAR__2540[7:0] ;
assign n769____DOLLAR__2548 =  ( $signed( n733____DOLLAR__2422 ) >>> ( 8'd4 ))  ;
assign n770____DOLLAR__2551 =  ( n768____DOLLAR__2549 ) ^ ( n769____DOLLAR__2548 )  ;
assign n771____DOLLAR__2552 =  ( n770____DOLLAR__2551 ) & ( 8'd15 )  ;
assign n772____DOLLAR__2657 =  ( n771____DOLLAR__2552 ) == ( 8'd15 )  ;
assign n773____DOLLAR__2650 =  ( n771____DOLLAR__2552 ) == ( 8'd14 )  ;
assign n774____DOLLAR__2643 =  ( n771____DOLLAR__2552 ) == ( 8'd13 )  ;
assign n775____DOLLAR__2636 =  ( n771____DOLLAR__2552 ) == ( 8'd12 )  ;
assign n776____DOLLAR__2629 =  ( n771____DOLLAR__2552 ) == ( 8'd11 )  ;
assign n777____DOLLAR__2622 =  ( n771____DOLLAR__2552 ) == ( 8'd10 )  ;
assign n778____DOLLAR__2615 =  ( n771____DOLLAR__2552 ) == ( 8'd9 )  ;
assign n779____DOLLAR__2608 =  ( n771____DOLLAR__2552 ) == ( 8'd8 )  ;
assign n780____DOLLAR__2601 =  ( n771____DOLLAR__2552 ) == ( 8'd7 )  ;
assign n781____DOLLAR__2594 =  ( n771____DOLLAR__2552 ) == ( 8'd6 )  ;
assign n782____DOLLAR__2587 =  ( n771____DOLLAR__2552 ) == ( 8'd5 )  ;
assign n783____DOLLAR__2580 =  ( n771____DOLLAR__2552 ) == ( 8'd4 )  ;
assign n784____DOLLAR__2573 =  ( n771____DOLLAR__2552 ) == ( 8'd3 )  ;
assign n785____DOLLAR__2566 =  ( n771____DOLLAR__2552 ) == ( 8'd2 )  ;
assign n786____DOLLAR__2559 =  ( n771____DOLLAR__2552 ) == ( 8'd1 )  ;
assign n787____DOLLAR__2561 =  ( n786____DOLLAR__2559 ) ? ( 32'd498536548 ) : ( 32'd0 ) ;
assign n788____DOLLAR__2568 =  ( n785____DOLLAR__2566 ) ? ( 32'd997073096 ) : ( n787____DOLLAR__2561 ) ;
assign n789____DOLLAR__2575 =  ( n784____DOLLAR__2573 ) ? ( 32'd651767980 ) : ( n788____DOLLAR__2568 ) ;
assign n790____DOLLAR__2582 =  ( n783____DOLLAR__2580 ) ? ( 32'd1994146192 ) : ( n789____DOLLAR__2575 ) ;
assign n791____DOLLAR__2589 =  ( n782____DOLLAR__2587 ) ? ( 32'd1802195444 ) : ( n790____DOLLAR__2582 ) ;
assign n792____DOLLAR__2596 =  ( n781____DOLLAR__2594 ) ? ( 32'd1303535960 ) : ( n791____DOLLAR__2589 ) ;
assign n793____DOLLAR__2603 =  ( n780____DOLLAR__2601 ) ? ( 32'd1342533948 ) : ( n792____DOLLAR__2596 ) ;
assign n794____DOLLAR__2610 =  ( n779____DOLLAR__2608 ) ? ( 32'd-306674912 ) : ( n793____DOLLAR__2603 ) ;
assign n795____DOLLAR__2617 =  ( n778____DOLLAR__2615 ) ? ( 32'd-267414716 ) : ( n794____DOLLAR__2610 ) ;
assign n796____DOLLAR__2624 =  ( n777____DOLLAR__2622 ) ? ( 32'd-690576408 ) : ( n795____DOLLAR__2617 ) ;
assign n797____DOLLAR__2631 =  ( n776____DOLLAR__2629 ) ? ( 32'd-882789492 ) : ( n796____DOLLAR__2624 ) ;
assign n798____DOLLAR__2638 =  ( n775____DOLLAR__2636 ) ? ( 32'd-1687895376 ) : ( n797____DOLLAR__2631 ) ;
assign n799____DOLLAR__2645 =  ( n774____DOLLAR__2643 ) ? ( 32'd-2032938284 ) : ( n798____DOLLAR__2638 ) ;
assign n800____DOLLAR__2652 =  ( n773____DOLLAR__2650 ) ? ( 32'd-1609899400 ) : ( n799____DOLLAR__2645 ) ;
assign n801____DOLLAR__2659 =  ( n772____DOLLAR__2657 ) ? ( 32'd-1111625188 ) : ( n800____DOLLAR__2652 ) ;
assign n802____DOLLAR__2543 =  ( $signed( n767____DOLLAR__2540 ) >>> ( 32'd4 ))  ;
assign n803____DOLLAR__2660 =  ( n801____DOLLAR__2659 ) ^ ( n802____DOLLAR__2543 )  ;
assign n804____DOLLAR__2665 =  ( n227____DOLLAR__2663 ) ? ( n803____DOLLAR__2660 ) : ( CRC_IN ) ;
always @(posedge clk) begin
   if(rst) begin
       TXFIFO_FULL <= TXFIFO_FULL_randinit ;
       TXFIFO_WUSED_QWD <= TXFIFO_WUSED_QWD_randinit ;
       TXFIFO_BUFF_RD_PTR <= TXFIFO_BUFF_RD_PTR_randinit ;
       TXFIFO_BUFF_WR_PTR <= TXFIFO_BUFF_WR_PTR_randinit ;
       TXFIFO_RD_OUTPUT <= TXFIFO_RD_OUTPUT_randinit ;
       TX_STATE <= TX_STATE_randinit ;
       TX_STATE_ENCAP <= TX_STATE_ENCAP_randinit ;
       TX_B2B_CNTR <= TX_B2B_CNTR_randinit ;
       TX_PACKET_BYTE_CNT <= TX_PACKET_BYTE_CNT_randinit ;
       TX_WCNT <= TX_WCNT_randinit ;
       XGMII_DOUT_REG <= XGMII_DOUT_REG_randinit ;
       XGMII_COUT_REG <= XGMII_COUT_REG_randinit ;
       TX_PKT_SENT <= TX_PKT_SENT_randinit ;
       TX_BYTE_SENT <= TX_BYTE_SENT_randinit ;
       CRC <= CRC_randinit ;
       CRC_DAT_IN <= CRC_DAT_IN_randinit ;
       CRC_IN <= CRC_IN_randinit ;
       TX_WCNT_INI <= TX_WCNT_INI_randinit ;
       TX_BUF <= TX_BUF_randinit ;
       __COUNTER_start__n4 <= 0;
   end
   else if(__START__ && __ILA_TX_FUNC_valid__) begin
       if ( __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ ) begin 
           __COUNTER_start__n4 <= 1; end
       else if( (__COUNTER_start__n4 >= 1 ) && ( __COUNTER_start__n4 < 255 )) begin
           __COUNTER_start__n4 <= __COUNTER_start__n4 + 1; end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           TXFIFO_FULL <= TXFIFO_FULL ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           TXFIFO_WUSED_QWD <= n7____DOLLAR__506 ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           TXFIFO_BUFF_RD_PTR <= n12____DOLLAR__498 ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           TXFIFO_BUFF_WR_PTR <= TXFIFO_BUFF_WR_PTR ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           TXFIFO_RD_OUTPUT <= n15____DOLLAR__483 ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           TX_STATE <= n17____DOLLAR__3171 ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           TX_STATE_ENCAP <= n19____DOLLAR__3178 ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           TX_B2B_CNTR <= n22____DOLLAR__3162 ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           TX_PACKET_BYTE_CNT <= TX_PACKET_BYTE_CNT ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           TX_WCNT <= n23____DOLLAR__3181 ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           XGMII_DOUT_REG <= n107____DOLLAR__3154 ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           XGMII_COUT_REG <= n143____DOLLAR__2867 ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           TX_PKT_SENT <= TX_PKT_SENT ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           TX_BYTE_SENT <= TX_BYTE_SENT ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           CRC <= n158____DOLLAR__2707 ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           CRC_DAT_IN <= n226____DOLLAR__746 ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           CRC_IN <= n804____DOLLAR__2665 ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           TX_WCNT_INI <= TX_WCNT_INI ;
       end
       if (__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__) begin
           TX_BUF <= TXFIFO_RD_OUTPUT ;
       end
   end
end
endmodule
