module TX_FUNC(
MODE_10G,
MODE_1G,
MODE_2P5G,
MODE_5G,
RESETN,
TX_DATA,
TX_WE,
__ILA_TX_FUNC_grant__,
clk,
rst,
__ILA_TX_FUNC_acc_decode__,
__ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__,
__ILA_TX_FUNC_decode_of_SET_B2B_CNTR_10G__,
__ILA_TX_FUNC_decode_of_WR_PKT_LASTONE_10G__,
__ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__,
__ILA_TX_FUNC_valid__,
TXFIFO_BUFF_data_n59,
TXFIFO_BUFF_data_n65,
TXFIFO_BUFF_data_n144,
TXFIFO_BUFF_addr_n58,
TXFIFO_BUFF_addr_n64,
TXFIFO_BUFF_addr_n143,
TXFIFO_FULL,
TXFIFO_WUSED_QWD,
TXFIFO_BUFF_RD_PTR,
TXFIFO_BUFF_WR_PTR,
TXFIFO_RD_OUTPUT,
TXFIFO_RD_EN,
TXFIFO_RD_EMPTY,
TX_STATE,
TX_STATE_ENCAP,
TX_B2B_CNTR,
TX_B2B_OK,
TX_PACKET_BYTE_CNT,
TX_WCNT,
XGMII_DOUT_REG,
XGMII_COUT_REG,
TX_PKT_SENT,
TX_BYTE_SENT,
CRC,
CRC_DAT_IN,
CRC_IN,
TX_WCNT_INI,
TX_BUF,
TX_FUNC_INSTR
);
input            MODE_10G;
input            MODE_1G;
input            MODE_2P5G;
input            MODE_5G;
input            RESETN;
input     [63:0] TX_DATA;
input            TX_WE;
input      [3:0] __ILA_TX_FUNC_grant__;
input            clk;
input            rst;
input     [63:0] TXFIFO_BUFF_data_n59;
input     [63:0] TXFIFO_BUFF_data_n65;
input     [63:0] TXFIFO_BUFF_data_n144;
output      [3:0] __ILA_TX_FUNC_acc_decode__;
output            __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__;
output            __ILA_TX_FUNC_decode_of_SET_B2B_CNTR_10G__;
output            __ILA_TX_FUNC_decode_of_WR_PKT_LASTONE_10G__;
output            __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__;
output            __ILA_TX_FUNC_valid__;
output      [4:0] TXFIFO_BUFF_addr_n58;
output      [4:0] TXFIFO_BUFF_addr_n64;
output      [4:0] TXFIFO_BUFF_addr_n143;
output reg            TXFIFO_FULL;
output reg     [12:0] TXFIFO_WUSED_QWD;
output reg      [4:0] TXFIFO_BUFF_RD_PTR;
output reg      [4:0] TXFIFO_BUFF_WR_PTR;
output reg     [63:0] TXFIFO_RD_OUTPUT;
output reg            TXFIFO_RD_EN;
output reg            TXFIFO_RD_EMPTY;
output reg      [4:0] TX_STATE;
output reg      [7:0] TX_STATE_ENCAP;
output reg      [5:0] TX_B2B_CNTR;
output reg            TX_B2B_OK;
output reg     [15:0] TX_PACKET_BYTE_CNT;
output reg     [15:0] TX_WCNT;
output reg     [63:0] XGMII_DOUT_REG;
output reg      [7:0] XGMII_COUT_REG;
output reg     [31:0] TX_PKT_SENT;
output reg     [31:0] TX_BYTE_SENT;
output reg     [31:0] CRC;
output reg     [63:0] CRC_DAT_IN;
output reg     [31:0] CRC_IN;
output reg     [15:0] TX_WCNT_INI;
output reg     [63:0] TX_BUF;
output reg      [2:0] TX_FUNC_INSTR;
wire            MODE_10G;
wire            MODE_1G;
wire            MODE_2P5G;
wire            MODE_5G;
wire            RESETN;
wire      [4:0] TXFIFO_BUFF_addr_n143;
wire      [4:0] TXFIFO_BUFF_addr_n58;
wire      [4:0] TXFIFO_BUFF_addr_n64;
wire     [63:0] TXFIFO_BUFF_data_n144;
wire     [63:0] TXFIFO_BUFF_data_n59;
wire     [63:0] TXFIFO_BUFF_data_n65;
wire     [63:0] TX_DATA;
wire            TX_WE;
wire      [3:0] __ILA_TX_FUNC_acc_decode__;
wire            __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__;
wire            __ILA_TX_FUNC_decode_of_SET_B2B_CNTR_10G__;
wire            __ILA_TX_FUNC_decode_of_WR_PKT_LASTONE_10G__;
wire            __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__;
wire      [3:0] __ILA_TX_FUNC_grant__;
wire            __ILA_TX_FUNC_valid__;
wire            clk;
wire            n0;
wire            n1;
wire            n10;
wire     [12:0] n100;
wire     [31:0] n1000;
wire     [31:0] n1001;
wire     [31:0] n1002;
wire     [31:0] n1003;
wire     [31:0] n1004;
wire     [31:0] n1005;
wire     [31:0] n1006;
wire     [31:0] n1007;
wire     [31:0] n1008;
wire     [31:0] n1009;
wire     [12:0] n101;
wire     [31:0] n1010;
wire     [31:0] n1011;
wire     [31:0] n1012;
wire     [31:0] n1013;
wire     [31:0] n1014;
wire      [7:0] n1015;
wire     [39:0] n1016;
wire     [63:0] n1017;
wire            n1018;
wire     [15:0] n1019;
wire     [15:0] n102;
wire     [47:0] n1020;
wire     [63:0] n1021;
wire            n1022;
wire     [23:0] n1023;
wire     [55:0] n1024;
wire     [63:0] n1025;
wire            n1026;
wire     [31:0] n1027;
wire     [63:0] n1028;
wire            n1029;
wire     [15:0] n103;
wire     [23:0] n1030;
wire     [39:0] n1031;
wire     [63:0] n1032;
wire            n1033;
wire     [15:0] n1034;
wire     [47:0] n1035;
wire     [63:0] n1036;
wire      [7:0] n1037;
wire     [55:0] n1038;
wire     [63:0] n1039;
wire     [15:0] n104;
wire     [63:0] n1040;
wire     [63:0] n1041;
wire     [63:0] n1042;
wire     [63:0] n1043;
wire     [63:0] n1044;
wire     [63:0] n1045;
wire     [63:0] n1046;
wire            n1047;
wire            n1048;
wire     [63:0] n1049;
wire     [15:0] n105;
wire            n1050;
wire     [63:0] n1051;
wire            n1052;
wire     [63:0] n1053;
wire            n1054;
wire     [63:0] n1055;
wire            n1056;
wire     [63:0] n1057;
wire            n1058;
wire     [55:0] n1059;
wire     [15:0] n106;
wire      [7:0] n1060;
wire     [63:0] n1061;
wire            n1062;
wire     [47:0] n1063;
wire     [15:0] n1064;
wire     [63:0] n1065;
wire     [39:0] n1066;
wire     [23:0] n1067;
wire     [63:0] n1068;
wire     [63:0] n1069;
wire     [31:0] n107;
wire     [63:0] n1070;
wire     [63:0] n1071;
wire     [63:0] n1072;
wire     [63:0] n1073;
wire     [63:0] n1074;
wire     [63:0] n1075;
wire     [63:0] n1076;
wire     [63:0] n1077;
wire     [63:0] n1078;
wire     [63:0] n1079;
wire     [63:0] n108;
wire            n1080;
wire            n1081;
wire            n1082;
wire            n1083;
wire            n1084;
wire            n1085;
wire            n1086;
wire            n1087;
wire            n1088;
wire            n1089;
wire     [47:0] n109;
wire            n1090;
wire            n1091;
wire            n1092;
wire            n1093;
wire            n1094;
wire      [7:0] n1095;
wire      [7:0] n1096;
wire      [7:0] n1097;
wire      [7:0] n1098;
wire      [7:0] n1099;
wire            n11;
wire     [63:0] n110;
wire      [7:0] n1100;
wire      [7:0] n1101;
wire            n1102;
wire            n1103;
wire            n1104;
wire            n1105;
wire            n1106;
wire            n1107;
wire            n1108;
wire            n1109;
wire            n111;
wire      [7:0] n1110;
wire      [7:0] n1111;
wire      [7:0] n1112;
wire      [7:0] n1113;
wire      [7:0] n1114;
wire      [7:0] n1115;
wire      [7:0] n1116;
wire      [7:0] n1117;
wire      [7:0] n1118;
wire      [7:0] n1119;
wire            n112;
wire     [31:0] n1120;
wire     [31:0] n1121;
wire     [31:0] n1122;
wire      [2:0] n1123;
wire            n1124;
wire            n1125;
wire            n1126;
wire     [31:0] n1127;
wire            n1128;
wire            n1129;
wire            n113;
wire     [31:0] n1130;
wire            n1131;
wire            n1132;
wire     [31:0] n1133;
wire     [31:0] n1134;
wire     [31:0] n1135;
wire     [31:0] n1136;
wire     [31:0] n1137;
wire     [31:0] n1138;
wire     [31:0] n1139;
wire            n114;
wire            n1140;
wire            n1141;
wire            n1142;
wire      [7:0] n1143;
wire     [55:0] n1144;
wire     [63:0] n1145;
wire            n1146;
wire     [15:0] n1147;
wire     [47:0] n1148;
wire     [63:0] n1149;
wire            n115;
wire            n1150;
wire     [23:0] n1151;
wire     [39:0] n1152;
wire     [63:0] n1153;
wire            n1154;
wire     [31:0] n1155;
wire     [63:0] n1156;
wire            n1157;
wire     [39:0] n1158;
wire     [63:0] n1159;
wire      [4:0] n116;
wire            n1160;
wire     [47:0] n1161;
wire     [63:0] n1162;
wire     [55:0] n1163;
wire     [63:0] n1164;
wire     [63:0] n1165;
wire     [63:0] n1166;
wire     [63:0] n1167;
wire     [63:0] n1168;
wire     [63:0] n1169;
wire      [4:0] n117;
wire     [63:0] n1170;
wire     [63:0] n1171;
wire            n1172;
wire            n1173;
wire      [7:0] n1174;
wire     [55:0] n1175;
wire     [63:0] n1176;
wire            n1177;
wire     [15:0] n1178;
wire     [47:0] n1179;
wire      [4:0] n118;
wire     [63:0] n1180;
wire            n1181;
wire     [23:0] n1182;
wire     [39:0] n1183;
wire     [63:0] n1184;
wire            n1185;
wire     [31:0] n1186;
wire     [31:0] n1187;
wire     [63:0] n1188;
wire            n1189;
wire      [4:0] n119;
wire     [39:0] n1190;
wire     [23:0] n1191;
wire     [63:0] n1192;
wire            n1193;
wire     [47:0] n1194;
wire     [15:0] n1195;
wire     [63:0] n1196;
wire     [55:0] n1197;
wire      [7:0] n1198;
wire     [63:0] n1199;
wire            n12;
wire            n120;
wire     [63:0] n1200;
wire     [63:0] n1201;
wire     [63:0] n1202;
wire     [63:0] n1203;
wire     [63:0] n1204;
wire     [63:0] n1205;
wire     [63:0] n1206;
wire     [63:0] n1207;
wire            n1208;
wire     [31:0] n1209;
wire            n121;
wire            n1210;
wire            n1211;
wire     [31:0] n1212;
wire            n1213;
wire     [31:0] n1214;
wire            n1215;
wire     [31:0] n1216;
wire            n1217;
wire     [31:0] n1218;
wire            n1219;
wire            n122;
wire     [31:0] n1220;
wire     [31:0] n1221;
wire     [31:0] n1222;
wire     [31:0] n1223;
wire     [31:0] n1224;
wire     [31:0] n1225;
wire     [31:0] n1226;
wire     [31:0] n1227;
wire     [31:0] n1228;
wire     [15:0] n1229;
wire            n123;
wire            n124;
wire            n125;
wire            n126;
wire            n127;
wire            n128;
wire            n129;
wire            n13;
wire      [4:0] n130;
wire      [4:0] n131;
wire      [4:0] n132;
wire      [4:0] n133;
wire            n134;
wire            n135;
wire            n136;
wire      [4:0] n137;
wire      [4:0] n138;
wire      [4:0] n139;
wire            n14;
wire      [4:0] n140;
wire      [4:0] n141;
wire      [4:0] n142;
wire     [63:0] n145;
wire            n146;
wire            n147;
wire            n148;
wire            n149;
wire            n15;
wire            n150;
wire            n151;
wire            n152;
wire      [2:0] n153;
wire            n154;
wire            n155;
wire            n156;
wire      [7:0] n157;
wire      [7:0] n158;
wire      [7:0] n159;
wire            n16;
wire      [7:0] n160;
wire            n161;
wire     [31:0] n162;
wire            n163;
wire     [31:0] n164;
wire            n165;
wire     [31:0] n166;
wire            n167;
wire     [31:0] n168;
wire            n169;
wire            n17;
wire     [31:0] n170;
wire            n171;
wire     [31:0] n172;
wire            n173;
wire     [31:0] n174;
wire            n175;
wire     [31:0] n176;
wire            n177;
wire     [31:0] n178;
wire            n179;
wire            n18;
wire     [31:0] n180;
wire            n181;
wire     [31:0] n182;
wire            n183;
wire     [31:0] n184;
wire            n185;
wire     [31:0] n186;
wire            n187;
wire     [31:0] n188;
wire            n189;
wire            n19;
wire     [31:0] n190;
wire     [31:0] n191;
wire     [31:0] n192;
wire     [31:0] n193;
wire     [31:0] n194;
wire     [31:0] n195;
wire     [31:0] n196;
wire     [31:0] n197;
wire     [31:0] n198;
wire     [31:0] n199;
wire            n2;
wire            n20;
wire     [31:0] n200;
wire     [31:0] n201;
wire     [31:0] n202;
wire     [31:0] n203;
wire     [31:0] n204;
wire     [31:0] n205;
wire     [31:0] n206;
wire     [31:0] n207;
wire     [31:0] n208;
wire      [7:0] n209;
wire            n21;
wire      [7:0] n210;
wire      [7:0] n211;
wire      [7:0] n212;
wire            n213;
wire     [31:0] n214;
wire            n215;
wire     [31:0] n216;
wire            n217;
wire     [31:0] n218;
wire            n219;
wire            n22;
wire     [31:0] n220;
wire            n221;
wire     [31:0] n222;
wire            n223;
wire     [31:0] n224;
wire            n225;
wire     [31:0] n226;
wire            n227;
wire     [31:0] n228;
wire            n229;
wire            n23;
wire     [31:0] n230;
wire            n231;
wire     [31:0] n232;
wire            n233;
wire     [31:0] n234;
wire            n235;
wire     [31:0] n236;
wire            n237;
wire     [31:0] n238;
wire            n239;
wire            n24;
wire     [31:0] n240;
wire            n241;
wire     [31:0] n242;
wire     [31:0] n243;
wire     [31:0] n244;
wire     [31:0] n245;
wire     [31:0] n246;
wire     [31:0] n247;
wire     [31:0] n248;
wire     [31:0] n249;
wire            n25;
wire     [31:0] n250;
wire     [31:0] n251;
wire     [31:0] n252;
wire     [31:0] n253;
wire     [31:0] n254;
wire     [31:0] n255;
wire     [31:0] n256;
wire     [31:0] n257;
wire     [31:0] n258;
wire     [31:0] n259;
wire            n26;
wire     [31:0] n260;
wire      [7:0] n261;
wire      [7:0] n262;
wire      [7:0] n263;
wire      [7:0] n264;
wire            n265;
wire     [31:0] n266;
wire            n267;
wire     [31:0] n268;
wire            n269;
wire            n27;
wire     [31:0] n270;
wire            n271;
wire     [31:0] n272;
wire            n273;
wire     [31:0] n274;
wire            n275;
wire     [31:0] n276;
wire            n277;
wire     [31:0] n278;
wire            n279;
wire            n28;
wire     [31:0] n280;
wire            n281;
wire     [31:0] n282;
wire            n283;
wire     [31:0] n284;
wire            n285;
wire     [31:0] n286;
wire            n287;
wire     [31:0] n288;
wire            n289;
wire            n29;
wire     [31:0] n290;
wire            n291;
wire     [31:0] n292;
wire            n293;
wire     [31:0] n294;
wire     [31:0] n295;
wire     [31:0] n296;
wire     [31:0] n297;
wire     [31:0] n298;
wire     [31:0] n299;
wire            n3;
wire            n30;
wire     [31:0] n300;
wire     [31:0] n301;
wire     [31:0] n302;
wire     [31:0] n303;
wire     [31:0] n304;
wire     [31:0] n305;
wire     [31:0] n306;
wire     [31:0] n307;
wire     [31:0] n308;
wire     [31:0] n309;
wire            n31;
wire     [31:0] n310;
wire     [31:0] n311;
wire     [31:0] n312;
wire      [7:0] n313;
wire      [7:0] n314;
wire      [7:0] n315;
wire      [7:0] n316;
wire            n317;
wire     [31:0] n318;
wire            n319;
wire            n32;
wire     [31:0] n320;
wire            n321;
wire     [31:0] n322;
wire            n323;
wire     [31:0] n324;
wire            n325;
wire     [31:0] n326;
wire            n327;
wire     [31:0] n328;
wire            n329;
wire            n33;
wire     [31:0] n330;
wire            n331;
wire     [31:0] n332;
wire            n333;
wire     [31:0] n334;
wire            n335;
wire     [31:0] n336;
wire            n337;
wire     [31:0] n338;
wire            n339;
wire            n34;
wire     [31:0] n340;
wire            n341;
wire     [31:0] n342;
wire            n343;
wire     [31:0] n344;
wire            n345;
wire     [31:0] n346;
wire     [31:0] n347;
wire     [31:0] n348;
wire     [31:0] n349;
wire            n35;
wire     [31:0] n350;
wire     [31:0] n351;
wire     [31:0] n352;
wire     [31:0] n353;
wire     [31:0] n354;
wire     [31:0] n355;
wire     [31:0] n356;
wire     [31:0] n357;
wire     [31:0] n358;
wire     [31:0] n359;
wire            n36;
wire     [31:0] n360;
wire     [31:0] n361;
wire     [31:0] n362;
wire     [31:0] n363;
wire     [31:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire            n369;
wire     [12:0] n37;
wire     [31:0] n370;
wire            n371;
wire     [31:0] n372;
wire            n373;
wire     [31:0] n374;
wire            n375;
wire     [31:0] n376;
wire            n377;
wire     [31:0] n378;
wire            n379;
wire     [12:0] n38;
wire     [31:0] n380;
wire            n381;
wire     [31:0] n382;
wire            n383;
wire     [31:0] n384;
wire            n385;
wire     [31:0] n386;
wire            n387;
wire     [31:0] n388;
wire            n389;
wire     [12:0] n39;
wire     [31:0] n390;
wire            n391;
wire     [31:0] n392;
wire            n393;
wire     [31:0] n394;
wire            n395;
wire     [31:0] n396;
wire            n397;
wire     [31:0] n398;
wire     [31:0] n399;
wire            n4;
wire            n40;
wire     [31:0] n400;
wire     [31:0] n401;
wire     [31:0] n402;
wire     [31:0] n403;
wire     [31:0] n404;
wire     [31:0] n405;
wire     [31:0] n406;
wire     [31:0] n407;
wire     [31:0] n408;
wire     [31:0] n409;
wire     [12:0] n41;
wire     [31:0] n410;
wire     [31:0] n411;
wire     [31:0] n412;
wire     [31:0] n413;
wire     [31:0] n414;
wire     [31:0] n415;
wire     [31:0] n416;
wire      [7:0] n417;
wire      [7:0] n418;
wire      [7:0] n419;
wire     [12:0] n42;
wire      [7:0] n420;
wire            n421;
wire     [31:0] n422;
wire            n423;
wire     [31:0] n424;
wire            n425;
wire     [31:0] n426;
wire            n427;
wire     [31:0] n428;
wire            n429;
wire            n43;
wire     [31:0] n430;
wire            n431;
wire     [31:0] n432;
wire            n433;
wire     [31:0] n434;
wire            n435;
wire     [31:0] n436;
wire            n437;
wire     [31:0] n438;
wire            n439;
wire            n44;
wire     [31:0] n440;
wire            n441;
wire     [31:0] n442;
wire            n443;
wire     [31:0] n444;
wire            n445;
wire     [31:0] n446;
wire            n447;
wire     [31:0] n448;
wire            n449;
wire      [4:0] n45;
wire     [31:0] n450;
wire     [31:0] n451;
wire     [31:0] n452;
wire     [31:0] n453;
wire     [31:0] n454;
wire     [31:0] n455;
wire     [31:0] n456;
wire     [31:0] n457;
wire     [31:0] n458;
wire     [31:0] n459;
wire      [4:0] n46;
wire     [31:0] n460;
wire     [31:0] n461;
wire     [31:0] n462;
wire     [31:0] n463;
wire     [31:0] n464;
wire     [31:0] n465;
wire     [31:0] n466;
wire     [31:0] n467;
wire     [31:0] n468;
wire      [7:0] n469;
wire      [4:0] n47;
wire      [7:0] n470;
wire      [7:0] n471;
wire      [7:0] n472;
wire            n473;
wire     [31:0] n474;
wire            n475;
wire     [31:0] n476;
wire            n477;
wire     [31:0] n478;
wire            n479;
wire            n48;
wire     [31:0] n480;
wire            n481;
wire     [31:0] n482;
wire            n483;
wire     [31:0] n484;
wire            n485;
wire     [31:0] n486;
wire            n487;
wire     [31:0] n488;
wire            n489;
wire      [4:0] n49;
wire     [31:0] n490;
wire            n491;
wire     [31:0] n492;
wire            n493;
wire     [31:0] n494;
wire            n495;
wire     [31:0] n496;
wire            n497;
wire     [31:0] n498;
wire            n499;
wire            n5;
wire      [4:0] n50;
wire     [31:0] n500;
wire            n501;
wire     [31:0] n502;
wire     [31:0] n503;
wire     [31:0] n504;
wire     [31:0] n505;
wire     [31:0] n506;
wire     [31:0] n507;
wire     [31:0] n508;
wire     [31:0] n509;
wire            n51;
wire     [31:0] n510;
wire     [31:0] n511;
wire     [31:0] n512;
wire     [31:0] n513;
wire     [31:0] n514;
wire     [31:0] n515;
wire     [31:0] n516;
wire     [31:0] n517;
wire     [31:0] n518;
wire     [31:0] n519;
wire            n52;
wire     [31:0] n520;
wire      [7:0] n521;
wire      [7:0] n522;
wire      [7:0] n523;
wire      [7:0] n524;
wire            n525;
wire     [31:0] n526;
wire            n527;
wire     [31:0] n528;
wire            n529;
wire      [4:0] n53;
wire     [31:0] n530;
wire            n531;
wire     [31:0] n532;
wire            n533;
wire     [31:0] n534;
wire            n535;
wire     [31:0] n536;
wire            n537;
wire     [31:0] n538;
wire            n539;
wire      [4:0] n54;
wire     [31:0] n540;
wire            n541;
wire     [31:0] n542;
wire            n543;
wire     [31:0] n544;
wire            n545;
wire     [31:0] n546;
wire            n547;
wire     [31:0] n548;
wire            n549;
wire      [4:0] n55;
wire     [31:0] n550;
wire            n551;
wire     [31:0] n552;
wire            n553;
wire     [31:0] n554;
wire     [31:0] n555;
wire     [31:0] n556;
wire     [31:0] n557;
wire     [31:0] n558;
wire     [31:0] n559;
wire            n56;
wire     [31:0] n560;
wire     [31:0] n561;
wire     [31:0] n562;
wire     [31:0] n563;
wire     [31:0] n564;
wire     [31:0] n565;
wire     [31:0] n566;
wire     [31:0] n567;
wire     [31:0] n568;
wire     [31:0] n569;
wire      [4:0] n57;
wire     [31:0] n570;
wire     [31:0] n571;
wire     [31:0] n572;
wire      [7:0] n573;
wire      [7:0] n574;
wire      [7:0] n575;
wire      [7:0] n576;
wire            n577;
wire     [31:0] n578;
wire            n579;
wire     [31:0] n580;
wire            n581;
wire     [31:0] n582;
wire            n583;
wire     [31:0] n584;
wire            n585;
wire     [31:0] n586;
wire            n587;
wire     [31:0] n588;
wire            n589;
wire     [31:0] n590;
wire            n591;
wire     [31:0] n592;
wire            n593;
wire     [31:0] n594;
wire            n595;
wire     [31:0] n596;
wire            n597;
wire     [31:0] n598;
wire            n599;
wire            n6;
wire     [63:0] n60;
wire     [31:0] n600;
wire            n601;
wire     [31:0] n602;
wire            n603;
wire     [31:0] n604;
wire            n605;
wire     [31:0] n606;
wire     [31:0] n607;
wire     [31:0] n608;
wire     [31:0] n609;
wire            n61;
wire     [31:0] n610;
wire     [31:0] n611;
wire     [31:0] n612;
wire     [31:0] n613;
wire     [31:0] n614;
wire     [31:0] n615;
wire     [31:0] n616;
wire     [31:0] n617;
wire     [31:0] n618;
wire     [31:0] n619;
wire            n62;
wire     [31:0] n620;
wire     [31:0] n621;
wire     [31:0] n622;
wire     [31:0] n623;
wire     [31:0] n624;
wire      [7:0] n625;
wire      [7:0] n626;
wire      [7:0] n627;
wire      [7:0] n628;
wire            n629;
wire      [4:0] n63;
wire     [31:0] n630;
wire            n631;
wire     [31:0] n632;
wire            n633;
wire     [31:0] n634;
wire            n635;
wire     [31:0] n636;
wire            n637;
wire     [31:0] n638;
wire            n639;
wire     [31:0] n640;
wire            n641;
wire     [31:0] n642;
wire            n643;
wire     [31:0] n644;
wire            n645;
wire     [31:0] n646;
wire            n647;
wire     [31:0] n648;
wire            n649;
wire     [31:0] n650;
wire            n651;
wire     [31:0] n652;
wire            n653;
wire     [31:0] n654;
wire            n655;
wire     [31:0] n656;
wire            n657;
wire     [31:0] n658;
wire     [31:0] n659;
wire     [63:0] n66;
wire     [31:0] n660;
wire     [31:0] n661;
wire     [31:0] n662;
wire     [31:0] n663;
wire     [31:0] n664;
wire     [31:0] n665;
wire     [31:0] n666;
wire     [31:0] n667;
wire     [31:0] n668;
wire     [31:0] n669;
wire     [63:0] n67;
wire     [31:0] n670;
wire     [31:0] n671;
wire     [31:0] n672;
wire     [31:0] n673;
wire     [31:0] n674;
wire     [31:0] n675;
wire     [31:0] n676;
wire      [7:0] n677;
wire      [7:0] n678;
wire      [7:0] n679;
wire            n68;
wire      [7:0] n680;
wire            n681;
wire     [31:0] n682;
wire            n683;
wire     [31:0] n684;
wire            n685;
wire     [31:0] n686;
wire            n687;
wire     [31:0] n688;
wire            n689;
wire            n69;
wire     [31:0] n690;
wire            n691;
wire     [31:0] n692;
wire            n693;
wire     [31:0] n694;
wire            n695;
wire     [31:0] n696;
wire            n697;
wire     [31:0] n698;
wire            n699;
wire            n7;
wire            n70;
wire     [31:0] n700;
wire            n701;
wire     [31:0] n702;
wire            n703;
wire     [31:0] n704;
wire            n705;
wire     [31:0] n706;
wire            n707;
wire     [31:0] n708;
wire            n709;
wire            n71;
wire     [31:0] n710;
wire     [31:0] n711;
wire     [31:0] n712;
wire     [31:0] n713;
wire     [31:0] n714;
wire     [31:0] n715;
wire     [31:0] n716;
wire     [31:0] n717;
wire     [31:0] n718;
wire     [31:0] n719;
wire            n72;
wire     [31:0] n720;
wire     [31:0] n721;
wire     [31:0] n722;
wire     [31:0] n723;
wire     [31:0] n724;
wire     [31:0] n725;
wire     [31:0] n726;
wire     [31:0] n727;
wire     [31:0] n728;
wire      [7:0] n729;
wire            n73;
wire      [7:0] n730;
wire      [7:0] n731;
wire      [7:0] n732;
wire            n733;
wire     [31:0] n734;
wire            n735;
wire     [31:0] n736;
wire            n737;
wire     [31:0] n738;
wire            n739;
wire            n74;
wire     [31:0] n740;
wire            n741;
wire     [31:0] n742;
wire            n743;
wire     [31:0] n744;
wire            n745;
wire     [31:0] n746;
wire            n747;
wire     [31:0] n748;
wire            n749;
wire            n75;
wire     [31:0] n750;
wire            n751;
wire     [31:0] n752;
wire            n753;
wire     [31:0] n754;
wire            n755;
wire     [31:0] n756;
wire            n757;
wire     [31:0] n758;
wire            n759;
wire            n76;
wire     [31:0] n760;
wire            n761;
wire     [31:0] n762;
wire     [31:0] n763;
wire     [31:0] n764;
wire     [31:0] n765;
wire     [31:0] n766;
wire     [31:0] n767;
wire     [31:0] n768;
wire     [31:0] n769;
wire            n77;
wire     [31:0] n770;
wire     [31:0] n771;
wire     [31:0] n772;
wire     [31:0] n773;
wire     [31:0] n774;
wire     [31:0] n775;
wire     [31:0] n776;
wire     [31:0] n777;
wire     [31:0] n778;
wire     [31:0] n779;
wire            n78;
wire     [31:0] n780;
wire      [7:0] n781;
wire      [7:0] n782;
wire      [7:0] n783;
wire      [7:0] n784;
wire            n785;
wire     [31:0] n786;
wire            n787;
wire     [31:0] n788;
wire            n789;
wire      [4:0] n79;
wire     [31:0] n790;
wire            n791;
wire     [31:0] n792;
wire            n793;
wire     [31:0] n794;
wire            n795;
wire     [31:0] n796;
wire            n797;
wire     [31:0] n798;
wire            n799;
wire            n8;
wire            n80;
wire     [31:0] n800;
wire            n801;
wire     [31:0] n802;
wire            n803;
wire     [31:0] n804;
wire            n805;
wire     [31:0] n806;
wire            n807;
wire     [31:0] n808;
wire            n809;
wire      [7:0] n81;
wire     [31:0] n810;
wire            n811;
wire     [31:0] n812;
wire            n813;
wire     [31:0] n814;
wire     [31:0] n815;
wire     [31:0] n816;
wire     [31:0] n817;
wire     [31:0] n818;
wire     [31:0] n819;
wire            n82;
wire     [31:0] n820;
wire     [31:0] n821;
wire     [31:0] n822;
wire     [31:0] n823;
wire     [31:0] n824;
wire     [31:0] n825;
wire     [31:0] n826;
wire     [31:0] n827;
wire     [31:0] n828;
wire     [31:0] n829;
wire      [5:0] n83;
wire     [31:0] n830;
wire     [31:0] n831;
wire     [31:0] n832;
wire      [7:0] n833;
wire      [7:0] n834;
wire      [7:0] n835;
wire      [7:0] n836;
wire            n837;
wire     [31:0] n838;
wire            n839;
wire      [5:0] n84;
wire     [31:0] n840;
wire            n841;
wire     [31:0] n842;
wire            n843;
wire     [31:0] n844;
wire            n845;
wire     [31:0] n846;
wire            n847;
wire     [31:0] n848;
wire            n849;
wire            n85;
wire     [31:0] n850;
wire            n851;
wire     [31:0] n852;
wire            n853;
wire     [31:0] n854;
wire            n855;
wire     [31:0] n856;
wire            n857;
wire     [31:0] n858;
wire            n859;
wire            n86;
wire     [31:0] n860;
wire            n861;
wire     [31:0] n862;
wire            n863;
wire     [31:0] n864;
wire            n865;
wire     [31:0] n866;
wire     [31:0] n867;
wire     [31:0] n868;
wire     [31:0] n869;
wire            n87;
wire     [31:0] n870;
wire     [31:0] n871;
wire     [31:0] n872;
wire     [31:0] n873;
wire     [31:0] n874;
wire     [31:0] n875;
wire     [31:0] n876;
wire     [31:0] n877;
wire     [31:0] n878;
wire     [31:0] n879;
wire      [5:0] n88;
wire     [31:0] n880;
wire     [31:0] n881;
wire     [31:0] n882;
wire     [31:0] n883;
wire     [31:0] n884;
wire      [7:0] n885;
wire      [7:0] n886;
wire      [7:0] n887;
wire      [7:0] n888;
wire            n889;
wire      [5:0] n89;
wire     [31:0] n890;
wire            n891;
wire     [31:0] n892;
wire            n893;
wire     [31:0] n894;
wire            n895;
wire     [31:0] n896;
wire            n897;
wire     [31:0] n898;
wire            n899;
wire            n9;
wire            n90;
wire     [31:0] n900;
wire            n901;
wire     [31:0] n902;
wire            n903;
wire     [31:0] n904;
wire            n905;
wire     [31:0] n906;
wire            n907;
wire     [31:0] n908;
wire            n909;
wire            n91;
wire     [31:0] n910;
wire            n911;
wire     [31:0] n912;
wire            n913;
wire     [31:0] n914;
wire            n915;
wire     [31:0] n916;
wire            n917;
wire     [31:0] n918;
wire     [31:0] n919;
wire            n92;
wire     [31:0] n920;
wire     [31:0] n921;
wire     [31:0] n922;
wire     [31:0] n923;
wire     [31:0] n924;
wire     [31:0] n925;
wire     [31:0] n926;
wire     [31:0] n927;
wire     [31:0] n928;
wire     [31:0] n929;
wire      [5:0] n93;
wire     [31:0] n930;
wire     [31:0] n931;
wire     [31:0] n932;
wire     [31:0] n933;
wire     [31:0] n934;
wire     [31:0] n935;
wire     [31:0] n936;
wire      [7:0] n937;
wire      [7:0] n938;
wire      [7:0] n939;
wire      [5:0] n94;
wire      [7:0] n940;
wire            n941;
wire     [31:0] n942;
wire            n943;
wire     [31:0] n944;
wire            n945;
wire     [31:0] n946;
wire            n947;
wire     [31:0] n948;
wire            n949;
wire            n95;
wire     [31:0] n950;
wire            n951;
wire     [31:0] n952;
wire            n953;
wire     [31:0] n954;
wire            n955;
wire     [31:0] n956;
wire            n957;
wire     [31:0] n958;
wire            n959;
wire            n96;
wire     [31:0] n960;
wire            n961;
wire     [31:0] n962;
wire            n963;
wire     [31:0] n964;
wire            n965;
wire     [31:0] n966;
wire            n967;
wire     [31:0] n968;
wire            n969;
wire     [15:0] n97;
wire     [31:0] n970;
wire     [31:0] n971;
wire     [31:0] n972;
wire     [31:0] n973;
wire     [31:0] n974;
wire     [31:0] n975;
wire     [31:0] n976;
wire     [31:0] n977;
wire     [31:0] n978;
wire     [31:0] n979;
wire      [2:0] n98;
wire     [31:0] n980;
wire     [31:0] n981;
wire     [31:0] n982;
wire     [31:0] n983;
wire     [31:0] n984;
wire     [31:0] n985;
wire     [31:0] n986;
wire     [31:0] n987;
wire     [31:0] n988;
wire     [31:0] n989;
wire            n99;
wire     [31:0] n990;
wire     [31:0] n991;
wire     [31:0] n992;
wire     [31:0] n993;
wire     [31:0] n994;
wire     [31:0] n995;
wire     [31:0] n996;
wire     [31:0] n997;
wire     [31:0] n998;
wire     [31:0] n999;
wire            rst;


assign __ILA_TX_FUNC_valid__ = 1'b1 ;
assign n0 =  ( MODE_10G ) == ( 1'b1 )  ;
assign n1 =  ( TX_STATE ) == ( 5'd1 )  ;
assign n2 =  ( n0 ) & (n1 )  ;
assign n3 =  ( TX_STATE_ENCAP ) == ( 8'd1 )  ;
assign n4 =  ( n2 ) & (n3 )  ;
assign n5 =  ( TX_B2B_CNTR ) == ( 6'd0 )  ;
assign n6 =  $signed( TX_B2B_CNTR ) > $signed( 6'd0 )  ;
assign n7 =  ( n5 ) | ( n6 )  ;
assign n8 =  ( n4 ) & (n7 )  ;
assign n9 =  ( TX_B2B_OK ) == ( 1'b0 )  ;
assign n10 =  ( n8 ) & (n9 )  ;
assign __ILA_TX_FUNC_decode_of_SET_B2B_CNTR_10G__ = n10 ;
assign __ILA_TX_FUNC_acc_decode__[0] = __ILA_TX_FUNC_decode_of_SET_B2B_CNTR_10G__ ;
assign n11 =  ( MODE_10G ) == ( 1'b1 )  ;
assign n12 =  ( TX_B2B_OK ) == ( 1'b1 )  ;
assign n13 =  ( n11 ) & (n12 )  ;
assign n14 =  ( TX_B2B_CNTR ) == ( 6'd0 )  ;
assign n15 =  ( n13 ) & (n14 )  ;
assign n16 =  ( TX_STATE ) == ( 5'd1 )  ;
assign n17 =  ( n15 ) & (n16 )  ;
assign n18 =  ( TX_STATE_ENCAP ) == ( 8'd1 )  ;
assign n19 =  ( n17 ) & (n18 )  ;
assign n20 =  ( TXFIFO_RD_EMPTY ) == ( 1'b0 )  ;
assign n21 =  ( n19 ) & (n20 )  ;
assign __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ = n21 ;
assign __ILA_TX_FUNC_acc_decode__[1] = __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ ;
assign n22 =  ( MODE_10G ) == ( 1'b1 )  ;
assign n23 =  ( TX_STATE ) == ( 5'd8 )  ;
assign n24 =  ( n22 ) & (n23 )  ;
assign n25 =  $signed( TX_WCNT ) > $signed( 16'd23 )  ;
assign n26 =  ( TXFIFO_RD_EMPTY ) == ( 1'b0 )  ;
assign n27 =  ( n25 ) & (n26 )  ;
assign n28 =  ( TX_WCNT ) == ( 16'd23 )  ;
assign n29 =  $signed( TX_WCNT ) < $signed( 16'd23 )  ;
assign n30 =  ( n28 ) | ( n29 )  ;
assign n31 =  ( n27 ) | ( n30 )  ;
assign n32 =  ( n24 ) & (n31 )  ;
assign __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ = n32 ;
assign __ILA_TX_FUNC_acc_decode__[2] = __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ ;
assign n33 =  ( MODE_10G ) == ( 1'b1 )  ;
assign n34 =  ( TX_STATE ) == ( 5'd16 )  ;
assign n35 =  ( n33 ) & (n34 )  ;
assign __ILA_TX_FUNC_decode_of_WR_PKT_LASTONE_10G__ = n35 ;
assign __ILA_TX_FUNC_acc_decode__[3] = __ILA_TX_FUNC_decode_of_WR_PKT_LASTONE_10G__ ;

// hand write assumptions for bug hunting
assign state_c1 = (TX_STATE == 5'd1) | (TX_STATE == 5'd8) | (TX_STATE == 5'd16);
assign state_c2 = (TX_STATE_ENCAP == 8'd1) | (TX_STATE_ENCAP == 8'd16);
assign state_c3 = ~(TX_STATE == 5'd1) | (TX_STATE_ENCAP == 8'd1);
assign state_c4 = ~(TX_STATE == 5'd8) | ((TX_STATE_ENCAP == 8'd1) | (TX_STATE_ENCAP == 8'd16));
assign state_c5 = ~(TX_STATE == 5'd16) | (TX_STATE_ENCAP == 8'd1);
assign wcnt_c1 = ~(TX_STATE == 5'd1) | (TX_WCNT == 16'd0);
assign b2b_not_neg = ( n5 ) | ( n6 );
assign b2b_ok_c1 = ~n6 | (TX_B2B_OK == 0);
assign no_empty = (TXFIFO_RD_EMPTY == 0);
assign not_empty_start = ~(TX_STATE == 5'd1) | (TXFIFO_RD_EMPTY == 0);
assign mode = (MODE_10G == 1);

assign instr_valid = __ILA_TX_FUNC_decode_of_SET_B2B_CNTR_10G__ | __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ | __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ | __ILA_TX_FUNC_decode_of_WR_PKT_LASTONE_10G__;


assign n36 =  ( TXFIFO_RD_EN ) == ( 1'b0 )  ;
assign n37 =  ( TXFIFO_WUSED_QWD ) - ( 13'd1 )  ;
assign n38 =  ( TXFIFO_WUSED_QWD ) - ( 13'd2 )  ;
assign n39 =  ( n36 ) ? ( n37 ) : ( n38 ) ;
assign n40 =  $signed( TX_WCNT ) > $signed( 16'd23 )  ;
assign n41 =  ( TXFIFO_WUSED_QWD ) - ( 13'd1 )  ;
assign n42 =  ( n40 ) ? ( n41 ) : ( TXFIFO_WUSED_QWD ) ;
assign n43 =  ( TXFIFO_RD_EN ) == ( 1'b0 )  ;
assign n44 =  ( TXFIFO_BUFF_RD_PTR ) == ( 5'd16 )  ;
assign n45 =  ( TXFIFO_BUFF_RD_PTR ) + ( 5'd1 )  ;
assign n46 =  ( n44 ) ? ( 5'd1 ) : ( n45 ) ;
assign n47 =  ( n43 ) ? ( TXFIFO_BUFF_RD_PTR ) : ( n46 ) ;
assign n48 =  ( n47 ) == ( 5'd16 )  ;
assign n49 =  ( n47 ) + ( 5'd1 )  ;
assign n50 =  ( n48 ) ? ( 5'd1 ) : ( n49 ) ;
assign n51 =  $signed( TX_WCNT ) > $signed( 16'd23 )  ;
assign n52 =  ( TXFIFO_BUFF_RD_PTR ) == ( 5'd16 )  ;
assign n53 =  ( TXFIFO_BUFF_RD_PTR ) + ( 5'd1 )  ;
assign n54 =  ( n52 ) ? ( 5'd1 ) : ( n53 ) ;
assign n55 =  ( n51 ) ? ( n54 ) : ( TXFIFO_BUFF_RD_PTR ) ;
assign n56 =  ( n47 ) == ( 5'd16 )  ;
assign n57 =  ( n56 ) ? ( 5'd0 ) : ( n47 ) ;
assign TXFIFO_BUFF_addr_n58 = n57 ;
assign n60 = TXFIFO_BUFF_data_n59 ;
assign n61 =  $signed( TX_WCNT ) > $signed( 16'd23 )  ;
assign n62 =  ( TXFIFO_BUFF_RD_PTR ) == ( 5'd16 )  ;
assign n63 =  ( n62 ) ? ( 5'd0 ) : ( TXFIFO_BUFF_RD_PTR ) ;
assign TXFIFO_BUFF_addr_n64 = n63 ;
assign n66 = TXFIFO_BUFF_data_n65 ;
assign n67 =  ( n61 ) ? ( n66 ) : ( TXFIFO_RD_OUTPUT ) ;
assign n68 =  ( TX_WE ) == ( 1'b0 )  ;
assign n69 =  ( TXFIFO_WUSED_QWD ) == ( 13'd1 )  ;
assign n70 =  ( n68 ) & (n69 )  ;
assign n71 =  ( n70 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n72 =  ( TX_WE ) == ( 1'b0 )  ;
assign n73 =  ( TXFIFO_WUSED_QWD ) == ( 13'd1 )  ;
assign n74 =  ( n72 ) & (n73 )  ;
assign n75 =  ( n74 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n76 =  ( TX_WCNT ) == ( 16'd0 )  ;
assign n77 =  $signed( TX_WCNT ) > $signed( 16'd0 )  ;
assign n78 =  ( n76 ) | ( n77 )  ;
assign n79 =  ( n78 ) ? ( 5'd8 ) : ( 5'd16 ) ;
assign n80 =  $signed( TX_WCNT ) < $signed( 16'd16 )  ;
assign n81 =  ( n80 ) ? ( 8'd1 ) : ( TX_STATE_ENCAP ) ;
assign n82 =  ( TX_B2B_CNTR ) == ( 6'd0 )  ;
assign n83 =  ( TX_B2B_CNTR ) - ( 6'd1 )  ;
assign n84 =  ( n82 ) ? ( TX_B2B_CNTR ) : ( n83 ) ;
assign n85 =  ( TX_STATE_ENCAP ) == ( 8'd1 )  ;
assign n86 =  $signed( TX_B2B_CNTR ) > $signed( 6'd0 )  ;
assign n87 =  ( n85 ) & (n86 )  ;
assign n88 =  ( TX_B2B_CNTR ) - ( 6'd1 )  ;
assign n89 =  ( n87 ) ? ( n88 ) : ( TX_B2B_CNTR ) ;
assign n90 =  ( TX_STATE_ENCAP ) == ( 8'd1 )  ;
assign n91 =  $signed( TX_B2B_CNTR ) > $signed( 6'd0 )  ;
assign n92 =  ( n90 ) & (n91 )  ;
assign n93 =  ( TX_B2B_CNTR ) - ( 6'd1 )  ;
assign n94 =  ( n92 ) ? ( n93 ) : ( TX_B2B_CNTR ) ;
assign n95 =  ( TX_B2B_CNTR ) == ( 6'd0 )  ;
assign n96 =  ( n95 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n97 = n60[15:0] ;
assign n98 = n97[2:0] ;
assign n99 =  ( n98 ) > ( 3'd0 )  ;
assign n100 = n97[15:3] ;
assign n101 =  ( n100 ) + ( 13'd1 )  ;
assign n102 =  { ( n101 ) , ( 3'd0 ) }  ;
assign n103 =  { ( n100 ) , ( 3'd0 ) }  ;
assign n104 =  ( n99 ) ? ( n102 ) : ( n103 ) ;
assign n105 =  ( n104 ) - ( 16'd1 )  ;
assign n106 =  ( TX_WCNT ) - ( 16'd8 )  ;
assign n107 =  { ( 16'd1799 ) , ( 16'd1799 ) }  ;
assign n108 =  { ( n107 ) , ( 32'd117901063 ) }  ;
assign n109 =  { ( 16'd21845 ) , ( 32'd1431655931 ) }  ;
assign n110 =  { ( 16'd54613 ) , ( n109 ) }  ;
assign n111 =  $signed( TX_WCNT ) > $signed( 16'd7 )  ;
assign n112 =  $signed( TX_WCNT ) > $signed( 16'd15 )  ;
assign n113 =  ( TXFIFO_BUFF_RD_PTR ) == ( 5'd3 )  ;
assign n114 =  ( TXFIFO_BUFF_RD_PTR ) > ( 5'd3 )  ;
assign n115 =  ( n113 ) | ( n114 )  ;
assign n116 =  ( TXFIFO_BUFF_RD_PTR ) - ( 5'd3 )  ;
assign n117 =  ( 5'd3 ) - ( TXFIFO_BUFF_RD_PTR )  ;
assign n118 =  ( 5'd16 ) - ( n117 )  ;
assign n119 =  ( n115 ) ? ( n116 ) : ( n118 ) ;
assign n120 =  ( TX_WCNT ) == ( 16'd8 )  ;
assign n121 =  $signed( TX_WCNT ) > $signed( 16'd8 )  ;
assign n122 =  ( n120 ) | ( n121 )  ;
assign n123 =  ( TX_WCNT ) == ( 16'd15 )  ;
assign n124 =  $signed( TX_WCNT ) < $signed( 16'd15 )  ;
assign n125 =  ( n123 ) | ( n124 )  ;
assign n126 =  ( n122 ) & (n125 )  ;
assign n127 =  ( TXFIFO_BUFF_RD_PTR ) == ( 5'd2 )  ;
assign n128 =  ( TXFIFO_BUFF_RD_PTR ) > ( 5'd2 )  ;
assign n129 =  ( n127 ) | ( n128 )  ;
assign n130 =  ( TXFIFO_BUFF_RD_PTR ) - ( 5'd2 )  ;
assign n131 =  ( 5'd2 ) - ( TXFIFO_BUFF_RD_PTR )  ;
assign n132 =  ( 5'd16 ) - ( n131 )  ;
assign n133 =  ( n129 ) ? ( n130 ) : ( n132 ) ;
assign n134 =  ( TXFIFO_BUFF_RD_PTR ) == ( 5'd1 )  ;
assign n135 =  ( TXFIFO_BUFF_RD_PTR ) > ( 5'd1 )  ;
assign n136 =  ( n134 ) | ( n135 )  ;
assign n137 =  ( TXFIFO_BUFF_RD_PTR ) - ( 5'd1 )  ;
assign n138 =  ( 5'd1 ) - ( TXFIFO_BUFF_RD_PTR )  ;
assign n139 =  ( 5'd16 ) - ( n138 )  ;
assign n140 =  ( n136 ) ? ( n137 ) : ( n139 ) ;
assign n141 =  ( n126 ) ? ( n133 ) : ( n140 ) ;
assign n142 =  ( n112 ) ? ( n119 ) : ( n141 ) ;
assign TXFIFO_BUFF_addr_n143 = n142 ;
assign n145 = TXFIFO_BUFF_data_n144 ;
assign n146 =  ( TX_WCNT ) == ( 16'd0 )  ;
assign n147 =  $signed( TX_WCNT ) > $signed( 16'd0 )  ;
assign n148 =  ( n146 ) | ( n147 )  ;
assign n149 =  ( TX_WCNT ) == ( 16'd7 )  ;
assign n150 =  $signed( TX_WCNT ) < $signed( 16'd7 )  ;
assign n151 =  ( n149 ) | ( n150 )  ;
assign n152 =  ( n148 ) & (n151 )  ;
assign n153 = TX_PACKET_BYTE_CNT[2:0] ;
assign n154 =  ( n153 ) == ( 3'd0 )  ;
assign n155 =  ( n153 ) == ( 3'd1 )  ;
assign n156 =  $signed( TX_WCNT ) > $signed( 16'd0 )  ;
assign n157 = CRC_IN[7:0] ;
assign n158 = CRC_DAT_IN[7:0] ;
assign n159 =  ( n157 ) ^ ( n158 )  ;
assign n160 =  ( n159 ) & ( 8'd15 )  ;
assign n161 =  ( n160 ) == ( 8'd15 )  ;
assign n162 =  { ( 16'd48573 ) , ( 16'd61980 ) }  ;
assign n163 =  ( n160 ) == ( 8'd14 )  ;
assign n164 =  { ( 16'd40970 ) , ( 16'd57976 ) }  ;
assign n165 =  ( n160 ) == ( 8'd13 )  ;
assign n166 =  { ( 16'd34515 ) , ( 16'd53972 ) }  ;
assign n167 =  ( n160 ) == ( 8'd12 )  ;
assign n168 =  { ( 16'd39780 ) , ( 16'd49840 ) }  ;
assign n169 =  ( n160 ) == ( 8'd11 )  ;
assign n170 =  { ( 16'd52065 ) , ( 16'd45964 ) }  ;
assign n171 =  ( n160 ) == ( 8'd10 )  ;
assign n172 =  { ( 16'd54998 ) , ( 16'd41960 ) }  ;
assign n173 =  ( n160 ) == ( 8'd9 )  ;
assign n174 =  { ( 16'd61455 ) , ( 16'd37700 ) }  ;
assign n175 =  ( n160 ) == ( 8'd8 )  ;
assign n176 =  { ( 16'd60856 ) , ( 16'd33568 ) }  ;
assign n177 =  ( n160 ) == ( 8'd7 )  ;
assign n178 =  { ( 16'd20485 ) , ( 16'd28988 ) }  ;
assign n179 =  ( n160 ) == ( 8'd6 )  ;
assign n180 =  { ( 16'd19890 ) , ( 16'd24920 ) }  ;
assign n181 =  ( n160 ) == ( 8'd5 )  ;
assign n182 =  { ( 16'd27499 ) , ( 16'd20980 ) }  ;
assign n183 =  ( n160 ) == ( 8'd4 )  ;
assign n184 =  { ( 16'd30428 ) , ( 16'd16784 ) }  ;
assign n185 =  ( n160 ) == ( 8'd3 )  ;
assign n186 =  { ( 16'd9945 ) , ( 16'd12460 ) }  ;
assign n187 =  ( n160 ) == ( 8'd2 )  ;
assign n188 =  { ( 16'd15214 ) , ( 16'd8392 ) }  ;
assign n189 =  ( n160 ) == ( 8'd1 )  ;
assign n190 =  { ( 16'd7607 ) , ( 16'd4196 ) }  ;
assign n191 =  { ( 16'd0 ) , ( 16'd0 ) }  ;
assign n192 =  ( n189 ) ? ( n190 ) : ( n191 ) ;
assign n193 =  ( n187 ) ? ( n188 ) : ( n192 ) ;
assign n194 =  ( n185 ) ? ( n186 ) : ( n193 ) ;
assign n195 =  ( n183 ) ? ( n184 ) : ( n194 ) ;
assign n196 =  ( n181 ) ? ( n182 ) : ( n195 ) ;
assign n197 =  ( n179 ) ? ( n180 ) : ( n196 ) ;
assign n198 =  ( n177 ) ? ( n178 ) : ( n197 ) ;
assign n199 =  ( n175 ) ? ( n176 ) : ( n198 ) ;
assign n200 =  ( n173 ) ? ( n174 ) : ( n199 ) ;
assign n201 =  ( n171 ) ? ( n172 ) : ( n200 ) ;
assign n202 =  ( n169 ) ? ( n170 ) : ( n201 ) ;
assign n203 =  ( n167 ) ? ( n168 ) : ( n202 ) ;
assign n204 =  ( n165 ) ? ( n166 ) : ( n203 ) ;
assign n205 =  ( n163 ) ? ( n164 ) : ( n204 ) ;
assign n206 =  ( n161 ) ? ( n162 ) : ( n205 ) ;
assign n207 =  ( ( CRC_IN ) >> ( 32'd4 ))  ;
assign n208 =  ( n206 ) ^ ( n207 )  ;
assign n209 = n208[7:0] ;
assign n210 =  ( ( n158 ) >> ( 8'd4 ))  ;
assign n211 =  ( n209 ) ^ ( n210 )  ;
assign n212 =  ( n211 ) & ( 8'd15 )  ;
assign n213 =  ( n212 ) == ( 8'd15 )  ;
assign n214 =  { ( 16'd48573 ) , ( 16'd61980 ) }  ;
assign n215 =  ( n212 ) == ( 8'd14 )  ;
assign n216 =  { ( 16'd40970 ) , ( 16'd57976 ) }  ;
assign n217 =  ( n212 ) == ( 8'd13 )  ;
assign n218 =  { ( 16'd34515 ) , ( 16'd53972 ) }  ;
assign n219 =  ( n212 ) == ( 8'd12 )  ;
assign n220 =  { ( 16'd39780 ) , ( 16'd49840 ) }  ;
assign n221 =  ( n212 ) == ( 8'd11 )  ;
assign n222 =  { ( 16'd52065 ) , ( 16'd45964 ) }  ;
assign n223 =  ( n212 ) == ( 8'd10 )  ;
assign n224 =  { ( 16'd54998 ) , ( 16'd41960 ) }  ;
assign n225 =  ( n212 ) == ( 8'd9 )  ;
assign n226 =  { ( 16'd61455 ) , ( 16'd37700 ) }  ;
assign n227 =  ( n212 ) == ( 8'd8 )  ;
assign n228 =  { ( 16'd60856 ) , ( 16'd33568 ) }  ;
assign n229 =  ( n212 ) == ( 8'd7 )  ;
assign n230 =  { ( 16'd20485 ) , ( 16'd28988 ) }  ;
assign n231 =  ( n212 ) == ( 8'd6 )  ;
assign n232 =  { ( 16'd19890 ) , ( 16'd24920 ) }  ;
assign n233 =  ( n212 ) == ( 8'd5 )  ;
assign n234 =  { ( 16'd27499 ) , ( 16'd20980 ) }  ;
assign n235 =  ( n212 ) == ( 8'd4 )  ;
assign n236 =  { ( 16'd30428 ) , ( 16'd16784 ) }  ;
assign n237 =  ( n212 ) == ( 8'd3 )  ;
assign n238 =  { ( 16'd9945 ) , ( 16'd12460 ) }  ;
assign n239 =  ( n212 ) == ( 8'd2 )  ;
assign n240 =  { ( 16'd15214 ) , ( 16'd8392 ) }  ;
assign n241 =  ( n212 ) == ( 8'd1 )  ;
assign n242 =  { ( 16'd7607 ) , ( 16'd4196 ) }  ;
assign n243 =  { ( 16'd0 ) , ( 16'd0 ) }  ;
assign n244 =  ( n241 ) ? ( n242 ) : ( n243 ) ;
assign n245 =  ( n239 ) ? ( n240 ) : ( n244 ) ;
assign n246 =  ( n237 ) ? ( n238 ) : ( n245 ) ;
assign n247 =  ( n235 ) ? ( n236 ) : ( n246 ) ;
assign n248 =  ( n233 ) ? ( n234 ) : ( n247 ) ;
assign n249 =  ( n231 ) ? ( n232 ) : ( n248 ) ;
assign n250 =  ( n229 ) ? ( n230 ) : ( n249 ) ;
assign n251 =  ( n227 ) ? ( n228 ) : ( n250 ) ;
assign n252 =  ( n225 ) ? ( n226 ) : ( n251 ) ;
assign n253 =  ( n223 ) ? ( n224 ) : ( n252 ) ;
assign n254 =  ( n221 ) ? ( n222 ) : ( n253 ) ;
assign n255 =  ( n219 ) ? ( n220 ) : ( n254 ) ;
assign n256 =  ( n217 ) ? ( n218 ) : ( n255 ) ;
assign n257 =  ( n215 ) ? ( n216 ) : ( n256 ) ;
assign n258 =  ( n213 ) ? ( n214 ) : ( n257 ) ;
assign n259 =  ( ( n208 ) >> ( 32'd4 ))  ;
assign n260 =  ( n258 ) ^ ( n259 )  ;
assign n261 = n260[7:0] ;
assign n262 = CRC_DAT_IN[15:8] ;
assign n263 =  ( n261 ) ^ ( n262 )  ;
assign n264 =  ( n263 ) & ( 8'd15 )  ;
assign n265 =  ( n264 ) == ( 8'd15 )  ;
assign n266 =  { ( 16'd48573 ) , ( 16'd61980 ) }  ;
assign n267 =  ( n264 ) == ( 8'd14 )  ;
assign n268 =  { ( 16'd40970 ) , ( 16'd57976 ) }  ;
assign n269 =  ( n264 ) == ( 8'd13 )  ;
assign n270 =  { ( 16'd34515 ) , ( 16'd53972 ) }  ;
assign n271 =  ( n264 ) == ( 8'd12 )  ;
assign n272 =  { ( 16'd39780 ) , ( 16'd49840 ) }  ;
assign n273 =  ( n264 ) == ( 8'd11 )  ;
assign n274 =  { ( 16'd52065 ) , ( 16'd45964 ) }  ;
assign n275 =  ( n264 ) == ( 8'd10 )  ;
assign n276 =  { ( 16'd54998 ) , ( 16'd41960 ) }  ;
assign n277 =  ( n264 ) == ( 8'd9 )  ;
assign n278 =  { ( 16'd61455 ) , ( 16'd37700 ) }  ;
assign n279 =  ( n264 ) == ( 8'd8 )  ;
assign n280 =  { ( 16'd60856 ) , ( 16'd33568 ) }  ;
assign n281 =  ( n264 ) == ( 8'd7 )  ;
assign n282 =  { ( 16'd20485 ) , ( 16'd28988 ) }  ;
assign n283 =  ( n264 ) == ( 8'd6 )  ;
assign n284 =  { ( 16'd19890 ) , ( 16'd24920 ) }  ;
assign n285 =  ( n264 ) == ( 8'd5 )  ;
assign n286 =  { ( 16'd27499 ) , ( 16'd20980 ) }  ;
assign n287 =  ( n264 ) == ( 8'd4 )  ;
assign n288 =  { ( 16'd30428 ) , ( 16'd16784 ) }  ;
assign n289 =  ( n264 ) == ( 8'd3 )  ;
assign n290 =  { ( 16'd9945 ) , ( 16'd12460 ) }  ;
assign n291 =  ( n264 ) == ( 8'd2 )  ;
assign n292 =  { ( 16'd15214 ) , ( 16'd8392 ) }  ;
assign n293 =  ( n264 ) == ( 8'd1 )  ;
assign n294 =  { ( 16'd7607 ) , ( 16'd4196 ) }  ;
assign n295 =  { ( 16'd0 ) , ( 16'd0 ) }  ;
assign n296 =  ( n293 ) ? ( n294 ) : ( n295 ) ;
assign n297 =  ( n291 ) ? ( n292 ) : ( n296 ) ;
assign n298 =  ( n289 ) ? ( n290 ) : ( n297 ) ;
assign n299 =  ( n287 ) ? ( n288 ) : ( n298 ) ;
assign n300 =  ( n285 ) ? ( n286 ) : ( n299 ) ;
assign n301 =  ( n283 ) ? ( n284 ) : ( n300 ) ;
assign n302 =  ( n281 ) ? ( n282 ) : ( n301 ) ;
assign n303 =  ( n279 ) ? ( n280 ) : ( n302 ) ;
assign n304 =  ( n277 ) ? ( n278 ) : ( n303 ) ;
assign n305 =  ( n275 ) ? ( n276 ) : ( n304 ) ;
assign n306 =  ( n273 ) ? ( n274 ) : ( n305 ) ;
assign n307 =  ( n271 ) ? ( n272 ) : ( n306 ) ;
assign n308 =  ( n269 ) ? ( n270 ) : ( n307 ) ;
assign n309 =  ( n267 ) ? ( n268 ) : ( n308 ) ;
assign n310 =  ( n265 ) ? ( n266 ) : ( n309 ) ;
assign n311 =  ( ( n260 ) >> ( 32'd4 ))  ;
assign n312 =  ( n310 ) ^ ( n311 )  ;
assign n313 = n312[7:0] ;
assign n314 =  ( ( n262 ) >> ( 8'd4 ))  ;
assign n315 =  ( n313 ) ^ ( n314 )  ;
assign n316 =  ( n315 ) & ( 8'd15 )  ;
assign n317 =  ( n316 ) == ( 8'd15 )  ;
assign n318 =  { ( 16'd48573 ) , ( 16'd61980 ) }  ;
assign n319 =  ( n316 ) == ( 8'd14 )  ;
assign n320 =  { ( 16'd40970 ) , ( 16'd57976 ) }  ;
assign n321 =  ( n316 ) == ( 8'd13 )  ;
assign n322 =  { ( 16'd34515 ) , ( 16'd53972 ) }  ;
assign n323 =  ( n316 ) == ( 8'd12 )  ;
assign n324 =  { ( 16'd39780 ) , ( 16'd49840 ) }  ;
assign n325 =  ( n316 ) == ( 8'd11 )  ;
assign n326 =  { ( 16'd52065 ) , ( 16'd45964 ) }  ;
assign n327 =  ( n316 ) == ( 8'd10 )  ;
assign n328 =  { ( 16'd54998 ) , ( 16'd41960 ) }  ;
assign n329 =  ( n316 ) == ( 8'd9 )  ;
assign n330 =  { ( 16'd61455 ) , ( 16'd37700 ) }  ;
assign n331 =  ( n316 ) == ( 8'd8 )  ;
assign n332 =  { ( 16'd60856 ) , ( 16'd33568 ) }  ;
assign n333 =  ( n316 ) == ( 8'd7 )  ;
assign n334 =  { ( 16'd20485 ) , ( 16'd28988 ) }  ;
assign n335 =  ( n316 ) == ( 8'd6 )  ;
assign n336 =  { ( 16'd19890 ) , ( 16'd24920 ) }  ;
assign n337 =  ( n316 ) == ( 8'd5 )  ;
assign n338 =  { ( 16'd27499 ) , ( 16'd20980 ) }  ;
assign n339 =  ( n316 ) == ( 8'd4 )  ;
assign n340 =  { ( 16'd30428 ) , ( 16'd16784 ) }  ;
assign n341 =  ( n316 ) == ( 8'd3 )  ;
assign n342 =  { ( 16'd9945 ) , ( 16'd12460 ) }  ;
assign n343 =  ( n316 ) == ( 8'd2 )  ;
assign n344 =  { ( 16'd15214 ) , ( 16'd8392 ) }  ;
assign n345 =  ( n316 ) == ( 8'd1 )  ;
assign n346 =  { ( 16'd7607 ) , ( 16'd4196 ) }  ;
assign n347 =  { ( 16'd0 ) , ( 16'd0 ) }  ;
assign n348 =  ( n345 ) ? ( n346 ) : ( n347 ) ;
assign n349 =  ( n343 ) ? ( n344 ) : ( n348 ) ;
assign n350 =  ( n341 ) ? ( n342 ) : ( n349 ) ;
assign n351 =  ( n339 ) ? ( n340 ) : ( n350 ) ;
assign n352 =  ( n337 ) ? ( n338 ) : ( n351 ) ;
assign n353 =  ( n335 ) ? ( n336 ) : ( n352 ) ;
assign n354 =  ( n333 ) ? ( n334 ) : ( n353 ) ;
assign n355 =  ( n331 ) ? ( n332 ) : ( n354 ) ;
assign n356 =  ( n329 ) ? ( n330 ) : ( n355 ) ;
assign n357 =  ( n327 ) ? ( n328 ) : ( n356 ) ;
assign n358 =  ( n325 ) ? ( n326 ) : ( n357 ) ;
assign n359 =  ( n323 ) ? ( n324 ) : ( n358 ) ;
assign n360 =  ( n321 ) ? ( n322 ) : ( n359 ) ;
assign n361 =  ( n319 ) ? ( n320 ) : ( n360 ) ;
assign n362 =  ( n317 ) ? ( n318 ) : ( n361 ) ;
assign n363 =  ( ( n312 ) >> ( 32'd4 ))  ;
assign n364 =  ( n362 ) ^ ( n363 )  ;
assign n365 = n364[7:0] ;
assign n366 = CRC_DAT_IN[23:16] ;
assign n367 =  ( n365 ) ^ ( n366 )  ;
assign n368 =  ( n367 ) & ( 8'd15 )  ;
assign n369 =  ( n368 ) == ( 8'd15 )  ;
assign n370 =  { ( 16'd48573 ) , ( 16'd61980 ) }  ;
assign n371 =  ( n368 ) == ( 8'd14 )  ;
assign n372 =  { ( 16'd40970 ) , ( 16'd57976 ) }  ;
assign n373 =  ( n368 ) == ( 8'd13 )  ;
assign n374 =  { ( 16'd34515 ) , ( 16'd53972 ) }  ;
assign n375 =  ( n368 ) == ( 8'd12 )  ;
assign n376 =  { ( 16'd39780 ) , ( 16'd49840 ) }  ;
assign n377 =  ( n368 ) == ( 8'd11 )  ;
assign n378 =  { ( 16'd52065 ) , ( 16'd45964 ) }  ;
assign n379 =  ( n368 ) == ( 8'd10 )  ;
assign n380 =  { ( 16'd54998 ) , ( 16'd41960 ) }  ;
assign n381 =  ( n368 ) == ( 8'd9 )  ;
assign n382 =  { ( 16'd61455 ) , ( 16'd37700 ) }  ;
assign n383 =  ( n368 ) == ( 8'd8 )  ;
assign n384 =  { ( 16'd60856 ) , ( 16'd33568 ) }  ;
assign n385 =  ( n368 ) == ( 8'd7 )  ;
assign n386 =  { ( 16'd20485 ) , ( 16'd28988 ) }  ;
assign n387 =  ( n368 ) == ( 8'd6 )  ;
assign n388 =  { ( 16'd19890 ) , ( 16'd24920 ) }  ;
assign n389 =  ( n368 ) == ( 8'd5 )  ;
assign n390 =  { ( 16'd27499 ) , ( 16'd20980 ) }  ;
assign n391 =  ( n368 ) == ( 8'd4 )  ;
assign n392 =  { ( 16'd30428 ) , ( 16'd16784 ) }  ;
assign n393 =  ( n368 ) == ( 8'd3 )  ;
assign n394 =  { ( 16'd9945 ) , ( 16'd12460 ) }  ;
assign n395 =  ( n368 ) == ( 8'd2 )  ;
assign n396 =  { ( 16'd15214 ) , ( 16'd8392 ) }  ;
assign n397 =  ( n368 ) == ( 8'd1 )  ;
assign n398 =  { ( 16'd7607 ) , ( 16'd4196 ) }  ;
assign n399 =  { ( 16'd0 ) , ( 16'd0 ) }  ;
assign n400 =  ( n397 ) ? ( n398 ) : ( n399 ) ;
assign n401 =  ( n395 ) ? ( n396 ) : ( n400 ) ;
assign n402 =  ( n393 ) ? ( n394 ) : ( n401 ) ;
assign n403 =  ( n391 ) ? ( n392 ) : ( n402 ) ;
assign n404 =  ( n389 ) ? ( n390 ) : ( n403 ) ;
assign n405 =  ( n387 ) ? ( n388 ) : ( n404 ) ;
assign n406 =  ( n385 ) ? ( n386 ) : ( n405 ) ;
assign n407 =  ( n383 ) ? ( n384 ) : ( n406 ) ;
assign n408 =  ( n381 ) ? ( n382 ) : ( n407 ) ;
assign n409 =  ( n379 ) ? ( n380 ) : ( n408 ) ;
assign n410 =  ( n377 ) ? ( n378 ) : ( n409 ) ;
assign n411 =  ( n375 ) ? ( n376 ) : ( n410 ) ;
assign n412 =  ( n373 ) ? ( n374 ) : ( n411 ) ;
assign n413 =  ( n371 ) ? ( n372 ) : ( n412 ) ;
assign n414 =  ( n369 ) ? ( n370 ) : ( n413 ) ;
assign n415 =  ( ( n364 ) >> ( 32'd4 ))  ;
assign n416 =  ( n414 ) ^ ( n415 )  ;
assign n417 = n416[7:0] ;
assign n418 =  ( ( n366 ) >> ( 8'd4 ))  ;
assign n419 =  ( n417 ) ^ ( n418 )  ;
assign n420 =  ( n419 ) & ( 8'd15 )  ;
assign n421 =  ( n420 ) == ( 8'd15 )  ;
assign n422 =  { ( 16'd48573 ) , ( 16'd61980 ) }  ;
assign n423 =  ( n420 ) == ( 8'd14 )  ;
assign n424 =  { ( 16'd40970 ) , ( 16'd57976 ) }  ;
assign n425 =  ( n420 ) == ( 8'd13 )  ;
assign n426 =  { ( 16'd34515 ) , ( 16'd53972 ) }  ;
assign n427 =  ( n420 ) == ( 8'd12 )  ;
assign n428 =  { ( 16'd39780 ) , ( 16'd49840 ) }  ;
assign n429 =  ( n420 ) == ( 8'd11 )  ;
assign n430 =  { ( 16'd52065 ) , ( 16'd45964 ) }  ;
assign n431 =  ( n420 ) == ( 8'd10 )  ;
assign n432 =  { ( 16'd54998 ) , ( 16'd41960 ) }  ;
assign n433 =  ( n420 ) == ( 8'd9 )  ;
assign n434 =  { ( 16'd61455 ) , ( 16'd37700 ) }  ;
assign n435 =  ( n420 ) == ( 8'd8 )  ;
assign n436 =  { ( 16'd60856 ) , ( 16'd33568 ) }  ;
assign n437 =  ( n420 ) == ( 8'd7 )  ;
assign n438 =  { ( 16'd20485 ) , ( 16'd28988 ) }  ;
assign n439 =  ( n420 ) == ( 8'd6 )  ;
assign n440 =  { ( 16'd19890 ) , ( 16'd24920 ) }  ;
assign n441 =  ( n420 ) == ( 8'd5 )  ;
assign n442 =  { ( 16'd27499 ) , ( 16'd20980 ) }  ;
assign n443 =  ( n420 ) == ( 8'd4 )  ;
assign n444 =  { ( 16'd30428 ) , ( 16'd16784 ) }  ;
assign n445 =  ( n420 ) == ( 8'd3 )  ;
assign n446 =  { ( 16'd9945 ) , ( 16'd12460 ) }  ;
assign n447 =  ( n420 ) == ( 8'd2 )  ;
assign n448 =  { ( 16'd15214 ) , ( 16'd8392 ) }  ;
assign n449 =  ( n420 ) == ( 8'd1 )  ;
assign n450 =  { ( 16'd7607 ) , ( 16'd4196 ) }  ;
assign n451 =  { ( 16'd0 ) , ( 16'd0 ) }  ;
assign n452 =  ( n449 ) ? ( n450 ) : ( n451 ) ;
assign n453 =  ( n447 ) ? ( n448 ) : ( n452 ) ;
assign n454 =  ( n445 ) ? ( n446 ) : ( n453 ) ;
assign n455 =  ( n443 ) ? ( n444 ) : ( n454 ) ;
assign n456 =  ( n441 ) ? ( n442 ) : ( n455 ) ;
assign n457 =  ( n439 ) ? ( n440 ) : ( n456 ) ;
assign n458 =  ( n437 ) ? ( n438 ) : ( n457 ) ;
assign n459 =  ( n435 ) ? ( n436 ) : ( n458 ) ;
assign n460 =  ( n433 ) ? ( n434 ) : ( n459 ) ;
assign n461 =  ( n431 ) ? ( n432 ) : ( n460 ) ;
assign n462 =  ( n429 ) ? ( n430 ) : ( n461 ) ;
assign n463 =  ( n427 ) ? ( n428 ) : ( n462 ) ;
assign n464 =  ( n425 ) ? ( n426 ) : ( n463 ) ;
assign n465 =  ( n423 ) ? ( n424 ) : ( n464 ) ;
assign n466 =  ( n421 ) ? ( n422 ) : ( n465 ) ;
assign n467 =  ( ( n416 ) >> ( 32'd4 ))  ;
assign n468 =  ( n466 ) ^ ( n467 )  ;
assign n469 = n468[7:0] ;
assign n470 = CRC_DAT_IN[31:24] ;
assign n471 =  ( n469 ) ^ ( n470 )  ;
assign n472 =  ( n471 ) & ( 8'd15 )  ;
assign n473 =  ( n472 ) == ( 8'd15 )  ;
assign n474 =  { ( 16'd48573 ) , ( 16'd61980 ) }  ;
assign n475 =  ( n472 ) == ( 8'd14 )  ;
assign n476 =  { ( 16'd40970 ) , ( 16'd57976 ) }  ;
assign n477 =  ( n472 ) == ( 8'd13 )  ;
assign n478 =  { ( 16'd34515 ) , ( 16'd53972 ) }  ;
assign n479 =  ( n472 ) == ( 8'd12 )  ;
assign n480 =  { ( 16'd39780 ) , ( 16'd49840 ) }  ;
assign n481 =  ( n472 ) == ( 8'd11 )  ;
assign n482 =  { ( 16'd52065 ) , ( 16'd45964 ) }  ;
assign n483 =  ( n472 ) == ( 8'd10 )  ;
assign n484 =  { ( 16'd54998 ) , ( 16'd41960 ) }  ;
assign n485 =  ( n472 ) == ( 8'd9 )  ;
assign n486 =  { ( 16'd61455 ) , ( 16'd37700 ) }  ;
assign n487 =  ( n472 ) == ( 8'd8 )  ;
assign n488 =  { ( 16'd60856 ) , ( 16'd33568 ) }  ;
assign n489 =  ( n472 ) == ( 8'd7 )  ;
assign n490 =  { ( 16'd20485 ) , ( 16'd28988 ) }  ;
assign n491 =  ( n472 ) == ( 8'd6 )  ;
assign n492 =  { ( 16'd19890 ) , ( 16'd24920 ) }  ;
assign n493 =  ( n472 ) == ( 8'd5 )  ;
assign n494 =  { ( 16'd27499 ) , ( 16'd20980 ) }  ;
assign n495 =  ( n472 ) == ( 8'd4 )  ;
assign n496 =  { ( 16'd30428 ) , ( 16'd16784 ) }  ;
assign n497 =  ( n472 ) == ( 8'd3 )  ;
assign n498 =  { ( 16'd9945 ) , ( 16'd12460 ) }  ;
assign n499 =  ( n472 ) == ( 8'd2 )  ;
assign n500 =  { ( 16'd15214 ) , ( 16'd8392 ) }  ;
assign n501 =  ( n472 ) == ( 8'd1 )  ;
assign n502 =  { ( 16'd7607 ) , ( 16'd4196 ) }  ;
assign n503 =  { ( 16'd0 ) , ( 16'd0 ) }  ;
assign n504 =  ( n501 ) ? ( n502 ) : ( n503 ) ;
assign n505 =  ( n499 ) ? ( n500 ) : ( n504 ) ;
assign n506 =  ( n497 ) ? ( n498 ) : ( n505 ) ;
assign n507 =  ( n495 ) ? ( n496 ) : ( n506 ) ;
assign n508 =  ( n493 ) ? ( n494 ) : ( n507 ) ;
assign n509 =  ( n491 ) ? ( n492 ) : ( n508 ) ;
assign n510 =  ( n489 ) ? ( n490 ) : ( n509 ) ;
assign n511 =  ( n487 ) ? ( n488 ) : ( n510 ) ;
assign n512 =  ( n485 ) ? ( n486 ) : ( n511 ) ;
assign n513 =  ( n483 ) ? ( n484 ) : ( n512 ) ;
assign n514 =  ( n481 ) ? ( n482 ) : ( n513 ) ;
assign n515 =  ( n479 ) ? ( n480 ) : ( n514 ) ;
assign n516 =  ( n477 ) ? ( n478 ) : ( n515 ) ;
assign n517 =  ( n475 ) ? ( n476 ) : ( n516 ) ;
assign n518 =  ( n473 ) ? ( n474 ) : ( n517 ) ;
assign n519 =  ( ( n468 ) >> ( 32'd4 ))  ;
assign n520 =  ( n518 ) ^ ( n519 )  ;
assign n521 = n520[7:0] ;
assign n522 =  ( ( n470 ) >> ( 8'd4 ))  ;
assign n523 =  ( n521 ) ^ ( n522 )  ;
assign n524 =  ( n523 ) & ( 8'd15 )  ;
assign n525 =  ( n524 ) == ( 8'd15 )  ;
assign n526 =  { ( 16'd48573 ) , ( 16'd61980 ) }  ;
assign n527 =  ( n524 ) == ( 8'd14 )  ;
assign n528 =  { ( 16'd40970 ) , ( 16'd57976 ) }  ;
assign n529 =  ( n524 ) == ( 8'd13 )  ;
assign n530 =  { ( 16'd34515 ) , ( 16'd53972 ) }  ;
assign n531 =  ( n524 ) == ( 8'd12 )  ;
assign n532 =  { ( 16'd39780 ) , ( 16'd49840 ) }  ;
assign n533 =  ( n524 ) == ( 8'd11 )  ;
assign n534 =  { ( 16'd52065 ) , ( 16'd45964 ) }  ;
assign n535 =  ( n524 ) == ( 8'd10 )  ;
assign n536 =  { ( 16'd54998 ) , ( 16'd41960 ) }  ;
assign n537 =  ( n524 ) == ( 8'd9 )  ;
assign n538 =  { ( 16'd61455 ) , ( 16'd37700 ) }  ;
assign n539 =  ( n524 ) == ( 8'd8 )  ;
assign n540 =  { ( 16'd60856 ) , ( 16'd33568 ) }  ;
assign n541 =  ( n524 ) == ( 8'd7 )  ;
assign n542 =  { ( 16'd20485 ) , ( 16'd28988 ) }  ;
assign n543 =  ( n524 ) == ( 8'd6 )  ;
assign n544 =  { ( 16'd19890 ) , ( 16'd24920 ) }  ;
assign n545 =  ( n524 ) == ( 8'd5 )  ;
assign n546 =  { ( 16'd27499 ) , ( 16'd20980 ) }  ;
assign n547 =  ( n524 ) == ( 8'd4 )  ;
assign n548 =  { ( 16'd30428 ) , ( 16'd16784 ) }  ;
assign n549 =  ( n524 ) == ( 8'd3 )  ;
assign n550 =  { ( 16'd9945 ) , ( 16'd12460 ) }  ;
assign n551 =  ( n524 ) == ( 8'd2 )  ;
assign n552 =  { ( 16'd15214 ) , ( 16'd8392 ) }  ;
assign n553 =  ( n524 ) == ( 8'd1 )  ;
assign n554 =  { ( 16'd7607 ) , ( 16'd4196 ) }  ;
assign n555 =  { ( 16'd0 ) , ( 16'd0 ) }  ;
assign n556 =  ( n553 ) ? ( n554 ) : ( n555 ) ;
assign n557 =  ( n551 ) ? ( n552 ) : ( n556 ) ;
assign n558 =  ( n549 ) ? ( n550 ) : ( n557 ) ;
assign n559 =  ( n547 ) ? ( n548 ) : ( n558 ) ;
assign n560 =  ( n545 ) ? ( n546 ) : ( n559 ) ;
assign n561 =  ( n543 ) ? ( n544 ) : ( n560 ) ;
assign n562 =  ( n541 ) ? ( n542 ) : ( n561 ) ;
assign n563 =  ( n539 ) ? ( n540 ) : ( n562 ) ;
assign n564 =  ( n537 ) ? ( n538 ) : ( n563 ) ;
assign n565 =  ( n535 ) ? ( n536 ) : ( n564 ) ;
assign n566 =  ( n533 ) ? ( n534 ) : ( n565 ) ;
assign n567 =  ( n531 ) ? ( n532 ) : ( n566 ) ;
assign n568 =  ( n529 ) ? ( n530 ) : ( n567 ) ;
assign n569 =  ( n527 ) ? ( n528 ) : ( n568 ) ;
assign n570 =  ( n525 ) ? ( n526 ) : ( n569 ) ;
assign n571 =  ( ( n520 ) >> ( 32'd4 ))  ;
assign n572 =  ( n570 ) ^ ( n571 )  ;
assign n573 = n572[7:0] ;
assign n574 = CRC_DAT_IN[39:32] ;
assign n575 =  ( n573 ) ^ ( n574 )  ;
assign n576 =  ( n575 ) & ( 8'd15 )  ;
assign n577 =  ( n576 ) == ( 8'd15 )  ;
assign n578 =  { ( 16'd48573 ) , ( 16'd61980 ) }  ;
assign n579 =  ( n576 ) == ( 8'd14 )  ;
assign n580 =  { ( 16'd40970 ) , ( 16'd57976 ) }  ;
assign n581 =  ( n576 ) == ( 8'd13 )  ;
assign n582 =  { ( 16'd34515 ) , ( 16'd53972 ) }  ;
assign n583 =  ( n576 ) == ( 8'd12 )  ;
assign n584 =  { ( 16'd39780 ) , ( 16'd49840 ) }  ;
assign n585 =  ( n576 ) == ( 8'd11 )  ;
assign n586 =  { ( 16'd52065 ) , ( 16'd45964 ) }  ;
assign n587 =  ( n576 ) == ( 8'd10 )  ;
assign n588 =  { ( 16'd54998 ) , ( 16'd41960 ) }  ;
assign n589 =  ( n576 ) == ( 8'd9 )  ;
assign n590 =  { ( 16'd61455 ) , ( 16'd37700 ) }  ;
assign n591 =  ( n576 ) == ( 8'd8 )  ;
assign n592 =  { ( 16'd60856 ) , ( 16'd33568 ) }  ;
assign n593 =  ( n576 ) == ( 8'd7 )  ;
assign n594 =  { ( 16'd20485 ) , ( 16'd28988 ) }  ;
assign n595 =  ( n576 ) == ( 8'd6 )  ;
assign n596 =  { ( 16'd19890 ) , ( 16'd24920 ) }  ;
assign n597 =  ( n576 ) == ( 8'd5 )  ;
assign n598 =  { ( 16'd27499 ) , ( 16'd20980 ) }  ;
assign n599 =  ( n576 ) == ( 8'd4 )  ;
assign n600 =  { ( 16'd30428 ) , ( 16'd16784 ) }  ;
assign n601 =  ( n576 ) == ( 8'd3 )  ;
assign n602 =  { ( 16'd9945 ) , ( 16'd12460 ) }  ;
assign n603 =  ( n576 ) == ( 8'd2 )  ;
assign n604 =  { ( 16'd15214 ) , ( 16'd8392 ) }  ;
assign n605 =  ( n576 ) == ( 8'd1 )  ;
assign n606 =  { ( 16'd7607 ) , ( 16'd4196 ) }  ;
assign n607 =  { ( 16'd0 ) , ( 16'd0 ) }  ;
assign n608 =  ( n605 ) ? ( n606 ) : ( n607 ) ;
assign n609 =  ( n603 ) ? ( n604 ) : ( n608 ) ;
assign n610 =  ( n601 ) ? ( n602 ) : ( n609 ) ;
assign n611 =  ( n599 ) ? ( n600 ) : ( n610 ) ;
assign n612 =  ( n597 ) ? ( n598 ) : ( n611 ) ;
assign n613 =  ( n595 ) ? ( n596 ) : ( n612 ) ;
assign n614 =  ( n593 ) ? ( n594 ) : ( n613 ) ;
assign n615 =  ( n591 ) ? ( n592 ) : ( n614 ) ;
assign n616 =  ( n589 ) ? ( n590 ) : ( n615 ) ;
assign n617 =  ( n587 ) ? ( n588 ) : ( n616 ) ;
assign n618 =  ( n585 ) ? ( n586 ) : ( n617 ) ;
assign n619 =  ( n583 ) ? ( n584 ) : ( n618 ) ;
assign n620 =  ( n581 ) ? ( n582 ) : ( n619 ) ;
assign n621 =  ( n579 ) ? ( n580 ) : ( n620 ) ;
assign n622 =  ( n577 ) ? ( n578 ) : ( n621 ) ;
assign n623 =  ( ( n572 ) >> ( 32'd4 ))  ;
assign n624 =  ( n622 ) ^ ( n623 )  ;
assign n625 = n624[7:0] ;
assign n626 =  ( ( n574 ) >> ( 8'd4 ))  ;
assign n627 =  ( n625 ) ^ ( n626 )  ;
assign n628 =  ( n627 ) & ( 8'd15 )  ;
assign n629 =  ( n628 ) == ( 8'd15 )  ;
assign n630 =  { ( 16'd48573 ) , ( 16'd61980 ) }  ;
assign n631 =  ( n628 ) == ( 8'd14 )  ;
assign n632 =  { ( 16'd40970 ) , ( 16'd57976 ) }  ;
assign n633 =  ( n628 ) == ( 8'd13 )  ;
assign n634 =  { ( 16'd34515 ) , ( 16'd53972 ) }  ;
assign n635 =  ( n628 ) == ( 8'd12 )  ;
assign n636 =  { ( 16'd39780 ) , ( 16'd49840 ) }  ;
assign n637 =  ( n628 ) == ( 8'd11 )  ;
assign n638 =  { ( 16'd52065 ) , ( 16'd45964 ) }  ;
assign n639 =  ( n628 ) == ( 8'd10 )  ;
assign n640 =  { ( 16'd54998 ) , ( 16'd41960 ) }  ;
assign n641 =  ( n628 ) == ( 8'd9 )  ;
assign n642 =  { ( 16'd61455 ) , ( 16'd37700 ) }  ;
assign n643 =  ( n628 ) == ( 8'd8 )  ;
assign n644 =  { ( 16'd60856 ) , ( 16'd33568 ) }  ;
assign n645 =  ( n628 ) == ( 8'd7 )  ;
assign n646 =  { ( 16'd20485 ) , ( 16'd28988 ) }  ;
assign n647 =  ( n628 ) == ( 8'd6 )  ;
assign n648 =  { ( 16'd19890 ) , ( 16'd24920 ) }  ;
assign n649 =  ( n628 ) == ( 8'd5 )  ;
assign n650 =  { ( 16'd27499 ) , ( 16'd20980 ) }  ;
assign n651 =  ( n628 ) == ( 8'd4 )  ;
assign n652 =  { ( 16'd30428 ) , ( 16'd16784 ) }  ;
assign n653 =  ( n628 ) == ( 8'd3 )  ;
assign n654 =  { ( 16'd9945 ) , ( 16'd12460 ) }  ;
assign n655 =  ( n628 ) == ( 8'd2 )  ;
assign n656 =  { ( 16'd15214 ) , ( 16'd8392 ) }  ;
assign n657 =  ( n628 ) == ( 8'd1 )  ;
assign n658 =  { ( 16'd7607 ) , ( 16'd4196 ) }  ;
assign n659 =  { ( 16'd0 ) , ( 16'd0 ) }  ;
assign n660 =  ( n657 ) ? ( n658 ) : ( n659 ) ;
assign n661 =  ( n655 ) ? ( n656 ) : ( n660 ) ;
assign n662 =  ( n653 ) ? ( n654 ) : ( n661 ) ;
assign n663 =  ( n651 ) ? ( n652 ) : ( n662 ) ;
assign n664 =  ( n649 ) ? ( n650 ) : ( n663 ) ;
assign n665 =  ( n647 ) ? ( n648 ) : ( n664 ) ;
assign n666 =  ( n645 ) ? ( n646 ) : ( n665 ) ;
assign n667 =  ( n643 ) ? ( n644 ) : ( n666 ) ;
assign n668 =  ( n641 ) ? ( n642 ) : ( n667 ) ;
assign n669 =  ( n639 ) ? ( n640 ) : ( n668 ) ;
assign n670 =  ( n637 ) ? ( n638 ) : ( n669 ) ;
assign n671 =  ( n635 ) ? ( n636 ) : ( n670 ) ;
assign n672 =  ( n633 ) ? ( n634 ) : ( n671 ) ;
assign n673 =  ( n631 ) ? ( n632 ) : ( n672 ) ;
assign n674 =  ( n629 ) ? ( n630 ) : ( n673 ) ;
assign n675 =  ( ( n624 ) >> ( 32'd4 ))  ;
assign n676 =  ( n674 ) ^ ( n675 )  ;
assign n677 = n676[7:0] ;
assign n678 = CRC_DAT_IN[47:40] ;
assign n679 =  ( n677 ) ^ ( n678 )  ;
assign n680 =  ( n679 ) & ( 8'd15 )  ;
assign n681 =  ( n680 ) == ( 8'd15 )  ;
assign n682 =  { ( 16'd48573 ) , ( 16'd61980 ) }  ;
assign n683 =  ( n680 ) == ( 8'd14 )  ;
assign n684 =  { ( 16'd40970 ) , ( 16'd57976 ) }  ;
assign n685 =  ( n680 ) == ( 8'd13 )  ;
assign n686 =  { ( 16'd34515 ) , ( 16'd53972 ) }  ;
assign n687 =  ( n680 ) == ( 8'd12 )  ;
assign n688 =  { ( 16'd39780 ) , ( 16'd49840 ) }  ;
assign n689 =  ( n680 ) == ( 8'd11 )  ;
assign n690 =  { ( 16'd52065 ) , ( 16'd45964 ) }  ;
assign n691 =  ( n680 ) == ( 8'd10 )  ;
assign n692 =  { ( 16'd54998 ) , ( 16'd41960 ) }  ;
assign n693 =  ( n680 ) == ( 8'd9 )  ;
assign n694 =  { ( 16'd61455 ) , ( 16'd37700 ) }  ;
assign n695 =  ( n680 ) == ( 8'd8 )  ;
assign n696 =  { ( 16'd60856 ) , ( 16'd33568 ) }  ;
assign n697 =  ( n680 ) == ( 8'd7 )  ;
assign n698 =  { ( 16'd20485 ) , ( 16'd28988 ) }  ;
assign n699 =  ( n680 ) == ( 8'd6 )  ;
assign n700 =  { ( 16'd19890 ) , ( 16'd24920 ) }  ;
assign n701 =  ( n680 ) == ( 8'd5 )  ;
assign n702 =  { ( 16'd27499 ) , ( 16'd20980 ) }  ;
assign n703 =  ( n680 ) == ( 8'd4 )  ;
assign n704 =  { ( 16'd30428 ) , ( 16'd16784 ) }  ;
assign n705 =  ( n680 ) == ( 8'd3 )  ;
assign n706 =  { ( 16'd9945 ) , ( 16'd12460 ) }  ;
assign n707 =  ( n680 ) == ( 8'd2 )  ;
assign n708 =  { ( 16'd15214 ) , ( 16'd8392 ) }  ;
assign n709 =  ( n680 ) == ( 8'd1 )  ;
assign n710 =  { ( 16'd7607 ) , ( 16'd4196 ) }  ;
assign n711 =  { ( 16'd0 ) , ( 16'd0 ) }  ;
assign n712 =  ( n709 ) ? ( n710 ) : ( n711 ) ;
assign n713 =  ( n707 ) ? ( n708 ) : ( n712 ) ;
assign n714 =  ( n705 ) ? ( n706 ) : ( n713 ) ;
assign n715 =  ( n703 ) ? ( n704 ) : ( n714 ) ;
assign n716 =  ( n701 ) ? ( n702 ) : ( n715 ) ;
assign n717 =  ( n699 ) ? ( n700 ) : ( n716 ) ;
assign n718 =  ( n697 ) ? ( n698 ) : ( n717 ) ;
assign n719 =  ( n695 ) ? ( n696 ) : ( n718 ) ;
assign n720 =  ( n693 ) ? ( n694 ) : ( n719 ) ;
assign n721 =  ( n691 ) ? ( n692 ) : ( n720 ) ;
assign n722 =  ( n689 ) ? ( n690 ) : ( n721 ) ;
assign n723 =  ( n687 ) ? ( n688 ) : ( n722 ) ;
assign n724 =  ( n685 ) ? ( n686 ) : ( n723 ) ;
assign n725 =  ( n683 ) ? ( n684 ) : ( n724 ) ;
assign n726 =  ( n681 ) ? ( n682 ) : ( n725 ) ;
assign n727 =  ( ( n676 ) >> ( 32'd4 ))  ;
assign n728 =  ( n726 ) ^ ( n727 )  ;
assign n729 = n728[7:0] ;
assign n730 =  ( ( n678 ) >> ( 8'd4 ))  ;
assign n731 =  ( n729 ) ^ ( n730 )  ;
assign n732 =  ( n731 ) & ( 8'd15 )  ;
assign n733 =  ( n732 ) == ( 8'd15 )  ;
assign n734 =  { ( 16'd48573 ) , ( 16'd61980 ) }  ;
assign n735 =  ( n732 ) == ( 8'd14 )  ;
assign n736 =  { ( 16'd40970 ) , ( 16'd57976 ) }  ;
assign n737 =  ( n732 ) == ( 8'd13 )  ;
assign n738 =  { ( 16'd34515 ) , ( 16'd53972 ) }  ;
assign n739 =  ( n732 ) == ( 8'd12 )  ;
assign n740 =  { ( 16'd39780 ) , ( 16'd49840 ) }  ;
assign n741 =  ( n732 ) == ( 8'd11 )  ;
assign n742 =  { ( 16'd52065 ) , ( 16'd45964 ) }  ;
assign n743 =  ( n732 ) == ( 8'd10 )  ;
assign n744 =  { ( 16'd54998 ) , ( 16'd41960 ) }  ;
assign n745 =  ( n732 ) == ( 8'd9 )  ;
assign n746 =  { ( 16'd61455 ) , ( 16'd37700 ) }  ;
assign n747 =  ( n732 ) == ( 8'd8 )  ;
assign n748 =  { ( 16'd60856 ) , ( 16'd33568 ) }  ;
assign n749 =  ( n732 ) == ( 8'd7 )  ;
assign n750 =  { ( 16'd20485 ) , ( 16'd28988 ) }  ;
assign n751 =  ( n732 ) == ( 8'd6 )  ;
assign n752 =  { ( 16'd19890 ) , ( 16'd24920 ) }  ;
assign n753 =  ( n732 ) == ( 8'd5 )  ;
assign n754 =  { ( 16'd27499 ) , ( 16'd20980 ) }  ;
assign n755 =  ( n732 ) == ( 8'd4 )  ;
assign n756 =  { ( 16'd30428 ) , ( 16'd16784 ) }  ;
assign n757 =  ( n732 ) == ( 8'd3 )  ;
assign n758 =  { ( 16'd9945 ) , ( 16'd12460 ) }  ;
assign n759 =  ( n732 ) == ( 8'd2 )  ;
assign n760 =  { ( 16'd15214 ) , ( 16'd8392 ) }  ;
assign n761 =  ( n732 ) == ( 8'd1 )  ;
assign n762 =  { ( 16'd7607 ) , ( 16'd4196 ) }  ;
assign n763 =  { ( 16'd0 ) , ( 16'd0 ) }  ;
assign n764 =  ( n761 ) ? ( n762 ) : ( n763 ) ;
assign n765 =  ( n759 ) ? ( n760 ) : ( n764 ) ;
assign n766 =  ( n757 ) ? ( n758 ) : ( n765 ) ;
assign n767 =  ( n755 ) ? ( n756 ) : ( n766 ) ;
assign n768 =  ( n753 ) ? ( n754 ) : ( n767 ) ;
assign n769 =  ( n751 ) ? ( n752 ) : ( n768 ) ;
assign n770 =  ( n749 ) ? ( n750 ) : ( n769 ) ;
assign n771 =  ( n747 ) ? ( n748 ) : ( n770 ) ;
assign n772 =  ( n745 ) ? ( n746 ) : ( n771 ) ;
assign n773 =  ( n743 ) ? ( n744 ) : ( n772 ) ;
assign n774 =  ( n741 ) ? ( n742 ) : ( n773 ) ;
assign n775 =  ( n739 ) ? ( n740 ) : ( n774 ) ;
assign n776 =  ( n737 ) ? ( n738 ) : ( n775 ) ;
assign n777 =  ( n735 ) ? ( n736 ) : ( n776 ) ;
assign n778 =  ( n733 ) ? ( n734 ) : ( n777 ) ;
assign n779 =  ( ( n728 ) >> ( 32'd4 ))  ;
assign n780 =  ( n778 ) ^ ( n779 )  ;
assign n781 = n780[7:0] ;
assign n782 = CRC_DAT_IN[55:48] ;
assign n783 =  ( n781 ) ^ ( n782 )  ;
assign n784 =  ( n783 ) & ( 8'd15 )  ;
assign n785 =  ( n784 ) == ( 8'd15 )  ;
assign n786 =  { ( 16'd48573 ) , ( 16'd61980 ) }  ;
assign n787 =  ( n784 ) == ( 8'd14 )  ;
assign n788 =  { ( 16'd40970 ) , ( 16'd57976 ) }  ;
assign n789 =  ( n784 ) == ( 8'd13 )  ;
assign n790 =  { ( 16'd34515 ) , ( 16'd53972 ) }  ;
assign n791 =  ( n784 ) == ( 8'd12 )  ;
assign n792 =  { ( 16'd39780 ) , ( 16'd49840 ) }  ;
assign n793 =  ( n784 ) == ( 8'd11 )  ;
assign n794 =  { ( 16'd52065 ) , ( 16'd45964 ) }  ;
assign n795 =  ( n784 ) == ( 8'd10 )  ;
assign n796 =  { ( 16'd54998 ) , ( 16'd41960 ) }  ;
assign n797 =  ( n784 ) == ( 8'd9 )  ;
assign n798 =  { ( 16'd61455 ) , ( 16'd37700 ) }  ;
assign n799 =  ( n784 ) == ( 8'd8 )  ;
assign n800 =  { ( 16'd60856 ) , ( 16'd33568 ) }  ;
assign n801 =  ( n784 ) == ( 8'd7 )  ;
assign n802 =  { ( 16'd20485 ) , ( 16'd28988 ) }  ;
assign n803 =  ( n784 ) == ( 8'd6 )  ;
assign n804 =  { ( 16'd19890 ) , ( 16'd24920 ) }  ;
assign n805 =  ( n784 ) == ( 8'd5 )  ;
assign n806 =  { ( 16'd27499 ) , ( 16'd20980 ) }  ;
assign n807 =  ( n784 ) == ( 8'd4 )  ;
assign n808 =  { ( 16'd30428 ) , ( 16'd16784 ) }  ;
assign n809 =  ( n784 ) == ( 8'd3 )  ;
assign n810 =  { ( 16'd9945 ) , ( 16'd12460 ) }  ;
assign n811 =  ( n784 ) == ( 8'd2 )  ;
assign n812 =  { ( 16'd15214 ) , ( 16'd8392 ) }  ;
assign n813 =  ( n784 ) == ( 8'd1 )  ;
assign n814 =  { ( 16'd7607 ) , ( 16'd4196 ) }  ;
assign n815 =  { ( 16'd0 ) , ( 16'd0 ) }  ;
assign n816 =  ( n813 ) ? ( n814 ) : ( n815 ) ;
assign n817 =  ( n811 ) ? ( n812 ) : ( n816 ) ;
assign n818 =  ( n809 ) ? ( n810 ) : ( n817 ) ;
assign n819 =  ( n807 ) ? ( n808 ) : ( n818 ) ;
assign n820 =  ( n805 ) ? ( n806 ) : ( n819 ) ;
assign n821 =  ( n803 ) ? ( n804 ) : ( n820 ) ;
assign n822 =  ( n801 ) ? ( n802 ) : ( n821 ) ;
assign n823 =  ( n799 ) ? ( n800 ) : ( n822 ) ;
assign n824 =  ( n797 ) ? ( n798 ) : ( n823 ) ;
assign n825 =  ( n795 ) ? ( n796 ) : ( n824 ) ;
assign n826 =  ( n793 ) ? ( n794 ) : ( n825 ) ;
assign n827 =  ( n791 ) ? ( n792 ) : ( n826 ) ;
assign n828 =  ( n789 ) ? ( n790 ) : ( n827 ) ;
assign n829 =  ( n787 ) ? ( n788 ) : ( n828 ) ;
assign n830 =  ( n785 ) ? ( n786 ) : ( n829 ) ;
assign n831 =  ( ( n780 ) >> ( 32'd4 ))  ;
assign n832 =  ( n830 ) ^ ( n831 )  ;
assign n833 = n832[7:0] ;
assign n834 =  ( ( n782 ) >> ( 8'd4 ))  ;
assign n835 =  ( n833 ) ^ ( n834 )  ;
assign n836 =  ( n835 ) & ( 8'd15 )  ;
assign n837 =  ( n836 ) == ( 8'd15 )  ;
assign n838 =  { ( 16'd48573 ) , ( 16'd61980 ) }  ;
assign n839 =  ( n836 ) == ( 8'd14 )  ;
assign n840 =  { ( 16'd40970 ) , ( 16'd57976 ) }  ;
assign n841 =  ( n836 ) == ( 8'd13 )  ;
assign n842 =  { ( 16'd34515 ) , ( 16'd53972 ) }  ;
assign n843 =  ( n836 ) == ( 8'd12 )  ;
assign n844 =  { ( 16'd39780 ) , ( 16'd49840 ) }  ;
assign n845 =  ( n836 ) == ( 8'd11 )  ;
assign n846 =  { ( 16'd52065 ) , ( 16'd45964 ) }  ;
assign n847 =  ( n836 ) == ( 8'd10 )  ;
assign n848 =  { ( 16'd54998 ) , ( 16'd41960 ) }  ;
assign n849 =  ( n836 ) == ( 8'd9 )  ;
assign n850 =  { ( 16'd61455 ) , ( 16'd37700 ) }  ;
assign n851 =  ( n836 ) == ( 8'd8 )  ;
assign n852 =  { ( 16'd60856 ) , ( 16'd33568 ) }  ;
assign n853 =  ( n836 ) == ( 8'd7 )  ;
assign n854 =  { ( 16'd20485 ) , ( 16'd28988 ) }  ;
assign n855 =  ( n836 ) == ( 8'd6 )  ;
assign n856 =  { ( 16'd19890 ) , ( 16'd24920 ) }  ;
assign n857 =  ( n836 ) == ( 8'd5 )  ;
assign n858 =  { ( 16'd27499 ) , ( 16'd20980 ) }  ;
assign n859 =  ( n836 ) == ( 8'd4 )  ;
assign n860 =  { ( 16'd30428 ) , ( 16'd16784 ) }  ;
assign n861 =  ( n836 ) == ( 8'd3 )  ;
assign n862 =  { ( 16'd9945 ) , ( 16'd12460 ) }  ;
assign n863 =  ( n836 ) == ( 8'd2 )  ;
assign n864 =  { ( 16'd15214 ) , ( 16'd8392 ) }  ;
assign n865 =  ( n836 ) == ( 8'd1 )  ;
assign n866 =  { ( 16'd7607 ) , ( 16'd4196 ) }  ;
assign n867 =  { ( 16'd0 ) , ( 16'd0 ) }  ;
assign n868 =  ( n865 ) ? ( n866 ) : ( n867 ) ;
assign n869 =  ( n863 ) ? ( n864 ) : ( n868 ) ;
assign n870 =  ( n861 ) ? ( n862 ) : ( n869 ) ;
assign n871 =  ( n859 ) ? ( n860 ) : ( n870 ) ;
assign n872 =  ( n857 ) ? ( n858 ) : ( n871 ) ;
assign n873 =  ( n855 ) ? ( n856 ) : ( n872 ) ;
assign n874 =  ( n853 ) ? ( n854 ) : ( n873 ) ;
assign n875 =  ( n851 ) ? ( n852 ) : ( n874 ) ;
assign n876 =  ( n849 ) ? ( n850 ) : ( n875 ) ;
assign n877 =  ( n847 ) ? ( n848 ) : ( n876 ) ;
assign n878 =  ( n845 ) ? ( n846 ) : ( n877 ) ;
assign n879 =  ( n843 ) ? ( n844 ) : ( n878 ) ;
assign n880 =  ( n841 ) ? ( n842 ) : ( n879 ) ;
assign n881 =  ( n839 ) ? ( n840 ) : ( n880 ) ;
assign n882 =  ( n837 ) ? ( n838 ) : ( n881 ) ;
assign n883 =  ( ( n832 ) >> ( 32'd4 ))  ;
assign n884 =  ( n882 ) ^ ( n883 )  ;
assign n885 = n884[7:0] ;
assign n886 = CRC_DAT_IN[63:56] ;
assign n887 =  ( n885 ) ^ ( n886 )  ;
assign n888 =  ( n887 ) & ( 8'd15 )  ;
assign n889 =  ( n888 ) == ( 8'd15 )  ;
assign n890 =  { ( 16'd48573 ) , ( 16'd61980 ) }  ;
assign n891 =  ( n888 ) == ( 8'd14 )  ;
assign n892 =  { ( 16'd40970 ) , ( 16'd57976 ) }  ;
assign n893 =  ( n888 ) == ( 8'd13 )  ;
assign n894 =  { ( 16'd34515 ) , ( 16'd53972 ) }  ;
assign n895 =  ( n888 ) == ( 8'd12 )  ;
assign n896 =  { ( 16'd39780 ) , ( 16'd49840 ) }  ;
assign n897 =  ( n888 ) == ( 8'd11 )  ;
assign n898 =  { ( 16'd52065 ) , ( 16'd45964 ) }  ;
assign n899 =  ( n888 ) == ( 8'd10 )  ;
assign n900 =  { ( 16'd54998 ) , ( 16'd41960 ) }  ;
assign n901 =  ( n888 ) == ( 8'd9 )  ;
assign n902 =  { ( 16'd61455 ) , ( 16'd37700 ) }  ;
assign n903 =  ( n888 ) == ( 8'd8 )  ;
assign n904 =  { ( 16'd60856 ) , ( 16'd33568 ) }  ;
assign n905 =  ( n888 ) == ( 8'd7 )  ;
assign n906 =  { ( 16'd20485 ) , ( 16'd28988 ) }  ;
assign n907 =  ( n888 ) == ( 8'd6 )  ;
assign n908 =  { ( 16'd19890 ) , ( 16'd24920 ) }  ;
assign n909 =  ( n888 ) == ( 8'd5 )  ;
assign n910 =  { ( 16'd27499 ) , ( 16'd20980 ) }  ;
assign n911 =  ( n888 ) == ( 8'd4 )  ;
assign n912 =  { ( 16'd30428 ) , ( 16'd16784 ) }  ;
assign n913 =  ( n888 ) == ( 8'd3 )  ;
assign n914 =  { ( 16'd9945 ) , ( 16'd12460 ) }  ;
assign n915 =  ( n888 ) == ( 8'd2 )  ;
assign n916 =  { ( 16'd15214 ) , ( 16'd8392 ) }  ;
assign n917 =  ( n888 ) == ( 8'd1 )  ;
assign n918 =  { ( 16'd7607 ) , ( 16'd4196 ) }  ;
assign n919 =  { ( 16'd0 ) , ( 16'd0 ) }  ;
assign n920 =  ( n917 ) ? ( n918 ) : ( n919 ) ;
assign n921 =  ( n915 ) ? ( n916 ) : ( n920 ) ;
assign n922 =  ( n913 ) ? ( n914 ) : ( n921 ) ;
assign n923 =  ( n911 ) ? ( n912 ) : ( n922 ) ;
assign n924 =  ( n909 ) ? ( n910 ) : ( n923 ) ;
assign n925 =  ( n907 ) ? ( n908 ) : ( n924 ) ;
assign n926 =  ( n905 ) ? ( n906 ) : ( n925 ) ;
assign n927 =  ( n903 ) ? ( n904 ) : ( n926 ) ;
assign n928 =  ( n901 ) ? ( n902 ) : ( n927 ) ;
assign n929 =  ( n899 ) ? ( n900 ) : ( n928 ) ;
assign n930 =  ( n897 ) ? ( n898 ) : ( n929 ) ;
assign n931 =  ( n895 ) ? ( n896 ) : ( n930 ) ;
assign n932 =  ( n893 ) ? ( n894 ) : ( n931 ) ;
assign n933 =  ( n891 ) ? ( n892 ) : ( n932 ) ;
assign n934 =  ( n889 ) ? ( n890 ) : ( n933 ) ;
assign n935 =  ( ( n884 ) >> ( 32'd4 ))  ;
assign n936 =  ( n934 ) ^ ( n935 )  ;
assign n937 = n936[7:0] ;
assign n938 =  ( ( n886 ) >> ( 8'd4 ))  ;
assign n939 =  ( n937 ) ^ ( n938 )  ;
assign n940 =  ( n939 ) & ( 8'd15 )  ;
assign n941 =  ( n940 ) == ( 8'd15 )  ;
assign n942 =  { ( 16'd48573 ) , ( 16'd61980 ) }  ;
assign n943 =  ( n940 ) == ( 8'd14 )  ;
assign n944 =  { ( 16'd40970 ) , ( 16'd57976 ) }  ;
assign n945 =  ( n940 ) == ( 8'd13 )  ;
assign n946 =  { ( 16'd34515 ) , ( 16'd53972 ) }  ;
assign n947 =  ( n940 ) == ( 8'd12 )  ;
assign n948 =  { ( 16'd39780 ) , ( 16'd49840 ) }  ;
assign n949 =  ( n940 ) == ( 8'd11 )  ;
assign n950 =  { ( 16'd52065 ) , ( 16'd45964 ) }  ;
assign n951 =  ( n940 ) == ( 8'd10 )  ;
assign n952 =  { ( 16'd54998 ) , ( 16'd41960 ) }  ;
assign n953 =  ( n940 ) == ( 8'd9 )  ;
assign n954 =  { ( 16'd61455 ) , ( 16'd37700 ) }  ;
assign n955 =  ( n940 ) == ( 8'd8 )  ;
assign n956 =  { ( 16'd60856 ) , ( 16'd33568 ) }  ;
assign n957 =  ( n940 ) == ( 8'd7 )  ;
assign n958 =  { ( 16'd20485 ) , ( 16'd28988 ) }  ;
assign n959 =  ( n940 ) == ( 8'd6 )  ;
assign n960 =  { ( 16'd19890 ) , ( 16'd24920 ) }  ;
assign n961 =  ( n940 ) == ( 8'd5 )  ;
assign n962 =  { ( 16'd27499 ) , ( 16'd20980 ) }  ;
assign n963 =  ( n940 ) == ( 8'd4 )  ;
assign n964 =  { ( 16'd30428 ) , ( 16'd16784 ) }  ;
assign n965 =  ( n940 ) == ( 8'd3 )  ;
assign n966 =  { ( 16'd9945 ) , ( 16'd12460 ) }  ;
assign n967 =  ( n940 ) == ( 8'd2 )  ;
assign n968 =  { ( 16'd15214 ) , ( 16'd8392 ) }  ;
assign n969 =  ( n940 ) == ( 8'd1 )  ;
assign n970 =  { ( 16'd7607 ) , ( 16'd4196 ) }  ;
assign n971 =  { ( 16'd0 ) , ( 16'd0 ) }  ;
assign n972 =  ( n969 ) ? ( n970 ) : ( n971 ) ;
assign n973 =  ( n967 ) ? ( n968 ) : ( n972 ) ;
assign n974 =  ( n965 ) ? ( n966 ) : ( n973 ) ;
assign n975 =  ( n963 ) ? ( n964 ) : ( n974 ) ;
assign n976 =  ( n961 ) ? ( n962 ) : ( n975 ) ;
assign n977 =  ( n959 ) ? ( n960 ) : ( n976 ) ;
assign n978 =  ( n957 ) ? ( n958 ) : ( n977 ) ;
assign n979 =  ( n955 ) ? ( n956 ) : ( n978 ) ;
assign n980 =  ( n953 ) ? ( n954 ) : ( n979 ) ;
assign n981 =  ( n951 ) ? ( n952 ) : ( n980 ) ;
assign n982 =  ( n949 ) ? ( n950 ) : ( n981 ) ;
assign n983 =  ( n947 ) ? ( n948 ) : ( n982 ) ;
assign n984 =  ( n945 ) ? ( n946 ) : ( n983 ) ;
assign n985 =  ( n943 ) ? ( n944 ) : ( n984 ) ;
assign n986 =  ( n941 ) ? ( n942 ) : ( n985 ) ;
assign n987 =  ( ( n936 ) >> ( 32'd4 ))  ;
assign n988 =  ( n986 ) ^ ( n987 )  ;
assign n989 =  ( n156 ) ? ( n988 ) : ( CRC_IN ) ;
assign n990 =  ( ( n989 ) >> ( 32'd24 ))  ;
assign n991 =  ( n990 ) & ( 32'd255 )  ;
assign n992 =  ( ( n989 ) >> ( 32'd8 ))  ;
assign n993 =  ( n992 ) & ( 32'd65280 )  ;
assign n994 =  ( n991 ) | ( n993 )  ;
assign n995 =  ( n989 ) << ( 32'd8 )  ;
assign n996 =  ( n995 ) & ( 32'd16711680 )  ;
assign n997 =  ( n994 ) | ( n996 )  ;
assign n998 =  ( n989 ) << ( 32'd24 )  ;
assign n999 =  { ( 16'd65280 ) , ( 16'd0 ) }  ;
assign n1000 =  ( n998 ) & ( n999 )  ;
assign n1001 =  ( n997 ) | ( n1000 )  ;
assign n1002 = ~ ( n1001 ) ;
assign n1003 =  ( ( n1002 ) >> ( 32'd24 ))  ;
assign n1004 =  ( n1003 ) & ( 32'd255 )  ;
assign n1005 =  ( ( n1002 ) >> ( 32'd8 ))  ;
assign n1006 =  ( n1005 ) & ( 32'd65280 )  ;
assign n1007 =  ( n1004 ) | ( n1006 )  ;
assign n1008 =  ( n1002 ) << ( 32'd8 )  ;
assign n1009 =  ( n1008 ) & ( 32'd16711680 )  ;
assign n1010 =  ( n1007 ) | ( n1009 )  ;
assign n1011 =  ( n1002 ) << ( 32'd24 )  ;
assign n1012 =  { ( 16'd65280 ) , ( 16'd0 ) }  ;
assign n1013 =  ( n1011 ) & ( n1012 )  ;
assign n1014 =  ( n1010 ) | ( n1013 )  ;
assign n1015 = n145[7:0] ;
assign n1016 =  { ( n1014 ) , ( n1015 ) }  ;
assign n1017 =  { ( 24'd460797 ) , ( n1016 ) }  ;
assign n1018 =  ( n153 ) == ( 3'd2 )  ;
assign n1019 = n145[15:0] ;
assign n1020 =  { ( n1014 ) , ( n1019 ) }  ;
assign n1021 =  { ( 16'd2045 ) , ( n1020 ) }  ;
assign n1022 =  ( n153 ) == ( 3'd3 )  ;
assign n1023 = n145[23:0] ;
assign n1024 =  { ( n1014 ) , ( n1023 ) }  ;
assign n1025 =  { ( 8'd253 ) , ( n1024 ) }  ;
assign n1026 =  ( n153 ) == ( 3'd4 )  ;
assign n1027 = n145[31:0] ;
assign n1028 =  { ( n1014 ) , ( n1027 ) }  ;
assign n1029 =  ( n153 ) == ( 3'd5 )  ;
assign n1030 = n1014[23:0] ;
assign n1031 = n145[39:0] ;
assign n1032 =  { ( n1030 ) , ( n1031 ) }  ;
assign n1033 =  ( n153 ) == ( 3'd6 )  ;
assign n1034 = n1014[15:0] ;
assign n1035 = n145[47:0] ;
assign n1036 =  { ( n1034 ) , ( n1035 ) }  ;
assign n1037 = n1014[7:0] ;
assign n1038 = n145[55:0] ;
assign n1039 =  { ( n1037 ) , ( n1038 ) }  ;
assign n1040 =  ( n1033 ) ? ( n1036 ) : ( n1039 ) ;
assign n1041 =  ( n1029 ) ? ( n1032 ) : ( n1040 ) ;
assign n1042 =  ( n1026 ) ? ( n1028 ) : ( n1041 ) ;
assign n1043 =  ( n1022 ) ? ( n1025 ) : ( n1042 ) ;
assign n1044 =  ( n1018 ) ? ( n1021 ) : ( n1043 ) ;
assign n1045 =  ( n155 ) ? ( n1017 ) : ( n1044 ) ;
assign n1046 =  ( n154 ) ? ( n145 ) : ( n1045 ) ;
assign n1047 =  $signed( TX_WCNT ) < $signed( 16'd0 )  ;
assign n1048 =  ( n153 ) == ( 3'd0 )  ;
assign n1049 =  { ( 32'd117901309 ) , ( n1014 ) }  ;
assign n1050 =  ( n153 ) == ( 3'd1 )  ;
assign n1051 =  { ( 32'd117901063 ) , ( 32'd117901063 ) }  ;
assign n1052 =  ( n153 ) == ( 3'd2 )  ;
assign n1053 =  { ( 32'd117901063 ) , ( 32'd117901063 ) }  ;
assign n1054 =  ( n153 ) == ( 3'd3 )  ;
assign n1055 =  { ( 32'd117901063 ) , ( 32'd117901063 ) }  ;
assign n1056 =  ( n153 ) == ( 3'd4 )  ;
assign n1057 =  { ( 32'd117901063 ) , ( 32'd117901309 ) }  ;
assign n1058 =  ( n153 ) == ( 3'd5 )  ;
assign n1059 =  { ( 32'd117901063 ) , ( 24'd460797 ) }  ;
assign n1060 = n1014[31:24] ;
assign n1061 =  { ( n1059 ) , ( n1060 ) }  ;
assign n1062 =  ( n153 ) == ( 3'd6 )  ;
assign n1063 =  { ( 32'd117901063 ) , ( 16'd2045 ) }  ;
assign n1064 = n1014[31:16] ;
assign n1065 =  { ( n1063 ) , ( n1064 ) }  ;
assign n1066 =  { ( 32'd117901063 ) , ( 8'd253 ) }  ;
assign n1067 = n1014[31:8] ;
assign n1068 =  { ( n1066 ) , ( n1067 ) }  ;
assign n1069 =  ( n1062 ) ? ( n1065 ) : ( n1068 ) ;
assign n1070 =  ( n1058 ) ? ( n1061 ) : ( n1069 ) ;
assign n1071 =  ( n1056 ) ? ( n1057 ) : ( n1070 ) ;
assign n1072 =  ( n1054 ) ? ( n1055 ) : ( n1071 ) ;
assign n1073 =  ( n1052 ) ? ( n1053 ) : ( n1072 ) ;
assign n1074 =  ( n1050 ) ? ( n1051 ) : ( n1073 ) ;
assign n1075 =  ( n1048 ) ? ( n1049 ) : ( n1074 ) ;
assign n1076 =  { ( 32'd117901063 ) , ( 32'd117901063 ) }  ;
assign n1077 =  ( n1047 ) ? ( n1075 ) : ( n1076 ) ;
assign n1078 =  ( n152 ) ? ( n1046 ) : ( n1077 ) ;
assign n1079 =  ( n111 ) ? ( n145 ) : ( n1078 ) ;
assign n1080 =  $signed( TX_WCNT ) > $signed( 16'd7 )  ;
assign n1081 =  ( TX_WCNT ) == ( 16'd0 )  ;
assign n1082 =  $signed( TX_WCNT ) > $signed( 16'd0 )  ;
assign n1083 =  ( n1081 ) | ( n1082 )  ;
assign n1084 =  ( TX_WCNT ) == ( 16'd7 )  ;
assign n1085 =  $signed( TX_WCNT ) < $signed( 16'd7 )  ;
assign n1086 =  ( n1084 ) | ( n1085 )  ;
assign n1087 =  ( n1083 ) & (n1086 )  ;
assign n1088 =  ( n153 ) == ( 3'd0 )  ;
assign n1089 =  ( n153 ) == ( 3'd1 )  ;
assign n1090 =  ( n153 ) == ( 3'd2 )  ;
assign n1091 =  ( n153 ) == ( 3'd3 )  ;
assign n1092 =  ( n153 ) == ( 3'd4 )  ;
assign n1093 =  ( n153 ) == ( 3'd5 )  ;
assign n1094 =  ( n153 ) == ( 3'd6 )  ;
assign n1095 =  ( n1094 ) ? ( 8'd0 ) : ( 8'd0 ) ;
assign n1096 =  ( n1093 ) ? ( 8'd0 ) : ( n1095 ) ;
assign n1097 =  ( n1092 ) ? ( 8'd0 ) : ( n1096 ) ;
assign n1098 =  ( n1091 ) ? ( 8'd128 ) : ( n1097 ) ;
assign n1099 =  ( n1090 ) ? ( 8'd192 ) : ( n1098 ) ;
assign n1100 =  ( n1089 ) ? ( 8'd224 ) : ( n1099 ) ;
assign n1101 =  ( n1088 ) ? ( 8'd0 ) : ( n1100 ) ;
assign n1102 =  $signed( TX_WCNT ) < $signed( 16'd0 )  ;
assign n1103 =  ( n153 ) == ( 3'd0 )  ;
assign n1104 =  ( n153 ) == ( 3'd1 )  ;
assign n1105 =  ( n153 ) == ( 3'd2 )  ;
assign n1106 =  ( n153 ) == ( 3'd3 )  ;
assign n1107 =  ( n153 ) == ( 3'd4 )  ;
assign n1108 =  ( n153 ) == ( 3'd5 )  ;
assign n1109 =  ( n153 ) == ( 3'd6 )  ;
assign n1110 =  ( n1109 ) ? ( 8'd252 ) : ( 8'd248 ) ;
assign n1111 =  ( n1108 ) ? ( 8'd254 ) : ( n1110 ) ;
assign n1112 =  ( n1107 ) ? ( 8'd255 ) : ( n1111 ) ;
assign n1113 =  ( n1106 ) ? ( 8'd255 ) : ( n1112 ) ;
assign n1114 =  ( n1105 ) ? ( 8'd255 ) : ( n1113 ) ;
assign n1115 =  ( n1104 ) ? ( 8'd255 ) : ( n1114 ) ;
assign n1116 =  ( n1103 ) ? ( 8'd240 ) : ( n1115 ) ;
assign n1117 =  ( n1102 ) ? ( n1116 ) : ( 8'd255 ) ;
assign n1118 =  ( n1087 ) ? ( n1101 ) : ( n1117 ) ;
assign n1119 =  ( n1080 ) ? ( 8'd0 ) : ( n1118 ) ;
assign n1120 =  ( TX_PKT_SENT ) + ( 32'd1 )  ;
assign n1121 =  { ( 16'd0 ) , ( TX_PACKET_BYTE_CNT ) }  ;
assign n1122 =  ( TX_BYTE_SENT ) + ( n1121 )  ;
assign n1123 = TX_PACKET_BYTE_CNT[2:0] ;
assign n1124 =  ( n1123 ) == ( 3'd0 )  ;
assign n1125 =  ( n1123 ) == ( 3'd1 )  ;
assign n1126 =  ( n1123 ) == ( 3'd2 )  ;
assign n1127 =  { ( 16'd59746 ) , ( 16'd45904 ) }  ;
assign n1128 =  ( n1123 ) == ( 3'd3 )  ;
assign n1129 =  ( n1123 ) == ( 3'd4 )  ;
assign n1130 =  { ( 16'd40202 ) , ( 16'd55661 ) }  ;
assign n1131 =  ( n1123 ) == ( 3'd5 )  ;
assign n1132 =  ( n1123 ) == ( 3'd6 )  ;
assign n1133 =  ( n1132 ) ? ( 32'd1868751717 ) : ( 32'd644901391 ) ;
assign n1134 =  ( n1131 ) ? ( 32'd2128204124 ) : ( n1133 ) ;
assign n1135 =  ( n1129 ) ? ( n1130 ) : ( n1134 ) ;
assign n1136 =  ( n1128 ) ? ( 32'd856065035 ) : ( n1135 ) ;
assign n1137 =  ( n1126 ) ? ( n1127 ) : ( n1136 ) ;
assign n1138 =  ( n1125 ) ? ( 32'd1453685177 ) : ( n1137 ) ;
assign n1139 =  ( n1124 ) ? ( 32'd0 ) : ( n1138 ) ;
assign n1140 =  ( TX_WCNT ) == ( TX_WCNT_INI )  ;
assign n1141 =  ( n153 ) == ( 3'd0 )  ;
assign n1142 =  ( n153 ) == ( 3'd1 )  ;
assign n1143 = n145[7:0] ;
assign n1144 =  { ( 32'd0 ) , ( 24'd0 ) }  ;
assign n1145 =  { ( n1143 ) , ( n1144 ) }  ;
assign n1146 =  ( n153 ) == ( 3'd2 )  ;
assign n1147 = n145[15:0] ;
assign n1148 =  { ( 32'd0 ) , ( 16'd0 ) }  ;
assign n1149 =  { ( n1147 ) , ( n1148 ) }  ;
assign n1150 =  ( n153 ) == ( 3'd3 )  ;
assign n1151 = n145[23:0] ;
assign n1152 =  { ( 32'd0 ) , ( 8'd0 ) }  ;
assign n1153 =  { ( n1151 ) , ( n1152 ) }  ;
assign n1154 =  ( n153 ) == ( 3'd4 )  ;
assign n1155 = n145[31:0] ;
assign n1156 =  { ( n1155 ) , ( 32'd0 ) }  ;
assign n1157 =  ( n153 ) == ( 3'd5 )  ;
assign n1158 = n145[39:0] ;
assign n1159 =  { ( n1158 ) , ( 24'd0 ) }  ;
assign n1160 =  ( n153 ) == ( 3'd6 )  ;
assign n1161 = n145[47:0] ;
assign n1162 =  { ( n1161 ) , ( 16'd0 ) }  ;
assign n1163 = n145[55:0] ;
assign n1164 =  { ( n1163 ) , ( 8'd0 ) }  ;
assign n1165 =  ( n1160 ) ? ( n1162 ) : ( n1164 ) ;
assign n1166 =  ( n1157 ) ? ( n1159 ) : ( n1165 ) ;
assign n1167 =  ( n1154 ) ? ( n1156 ) : ( n1166 ) ;
assign n1168 =  ( n1150 ) ? ( n1153 ) : ( n1167 ) ;
assign n1169 =  ( n1146 ) ? ( n1149 ) : ( n1168 ) ;
assign n1170 =  ( n1142 ) ? ( n1145 ) : ( n1169 ) ;
assign n1171 =  ( n1141 ) ? ( n145 ) : ( n1170 ) ;
assign n1172 =  ( n153 ) == ( 3'd0 )  ;
assign n1173 =  ( n153 ) == ( 3'd1 )  ;
assign n1174 = n145[7:0] ;
assign n1175 = TX_BUF[63:8] ;
assign n1176 =  { ( n1174 ) , ( n1175 ) }  ;
assign n1177 =  ( n153 ) == ( 3'd2 )  ;
assign n1178 = n145[15:0] ;
assign n1179 = TX_BUF[63:16] ;
assign n1180 =  { ( n1178 ) , ( n1179 ) }  ;
assign n1181 =  ( n153 ) == ( 3'd3 )  ;
assign n1182 = n145[23:0] ;
assign n1183 = TX_BUF[63:24] ;
assign n1184 =  { ( n1182 ) , ( n1183 ) }  ;
assign n1185 =  ( n153 ) == ( 3'd4 )  ;
assign n1186 = n145[31:0] ;
assign n1187 = TX_BUF[63:32] ;
assign n1188 =  { ( n1186 ) , ( n1187 ) }  ;
assign n1189 =  ( n153 ) == ( 3'd5 )  ;
assign n1190 = n145[39:0] ;
assign n1191 = TX_BUF[63:40] ;
assign n1192 =  { ( n1190 ) , ( n1191 ) }  ;
assign n1193 =  ( n153 ) == ( 3'd6 )  ;
assign n1194 = n145[47:0] ;
assign n1195 = TX_BUF[63:48] ;
assign n1196 =  { ( n1194 ) , ( n1195 ) }  ;
assign n1197 = n145[55:0] ;
assign n1198 = TX_BUF[63:56] ;
assign n1199 =  { ( n1197 ) , ( n1198 ) }  ;
assign n1200 =  ( n1193 ) ? ( n1196 ) : ( n1199 ) ;
assign n1201 =  ( n1189 ) ? ( n1192 ) : ( n1200 ) ;
assign n1202 =  ( n1185 ) ? ( n1188 ) : ( n1201 ) ;
assign n1203 =  ( n1181 ) ? ( n1184 ) : ( n1202 ) ;
assign n1204 =  ( n1177 ) ? ( n1180 ) : ( n1203 ) ;
assign n1205 =  ( n1173 ) ? ( n1176 ) : ( n1204 ) ;
assign n1206 =  ( n1172 ) ? ( n145 ) : ( n1205 ) ;
assign n1207 =  ( n1140 ) ? ( n1171 ) : ( n1206 ) ;
assign n1208 =  ( n1123 ) == ( 3'd0 )  ;
assign n1209 =  { ( 16'd65535 ) , ( 16'd65535 ) }  ;
assign n1210 =  ( n1123 ) == ( 3'd1 )  ;
assign n1211 =  ( n1123 ) == ( 3'd2 )  ;
assign n1212 =  { ( 16'd44876 ) , ( 16'd40214 ) }  ;
assign n1213 =  ( n1123 ) == ( 3'd3 )  ;
assign n1214 =  { ( 16'd62587 ) , ( 16'd63948 ) }  ;
assign n1215 =  ( n1123 ) == ( 3'd4 )  ;
assign n1216 =  { ( 16'd37414 ) , ( 16'd62818 ) }  ;
assign n1217 =  ( n1123 ) == ( 3'd5 )  ;
assign n1218 =  { ( 16'd41774 ) , ( 16'd9857 ) }  ;
assign n1219 =  ( n1123 ) == ( 3'd6 )  ;
assign n1220 =  { ( 16'd39452 ) , ( 16'd40336 ) }  ;
assign n1221 =  { ( 16'd61589 ) , ( 16'd36825 ) }  ;
assign n1222 =  ( n1219 ) ? ( n1220 ) : ( n1221 ) ;
assign n1223 =  ( n1217 ) ? ( n1218 ) : ( n1222 ) ;
assign n1224 =  ( n1215 ) ? ( n1216 ) : ( n1223 ) ;
assign n1225 =  ( n1213 ) ? ( n1214 ) : ( n1224 ) ;
assign n1226 =  ( n1211 ) ? ( n1212 ) : ( n1225 ) ;
assign n1227 =  ( n1210 ) ? ( 32'd1183210153 ) : ( n1226 ) ;
assign n1228 =  ( n1208 ) ? ( n1209 ) : ( n1227 ) ;
assign n1229 =  ( n104 ) - ( 16'd1 )  ;
always @(posedge clk) begin
   if(rst) begin
      TX_B2B_OK <= 1'b0;
      TX_B2B_CNTR <= 6'd6;
      TX_STATE <= 5'd1;
      TX_STATE_ENCAP <= 8'd1;
   end
   else if(__ILA_TX_FUNC_valid__) begin
       if ( __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ && __ILA_TX_FUNC_grant__[1] ) begin
           TXFIFO_WUSED_QWD <= n39;
       end else if ( __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ && __ILA_TX_FUNC_grant__[2] ) begin
           TXFIFO_WUSED_QWD <= n42;
       end
       if ( __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ && __ILA_TX_FUNC_grant__[1] ) begin
           TXFIFO_BUFF_RD_PTR <= n50;
       end else if ( __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ && __ILA_TX_FUNC_grant__[2] ) begin
           TXFIFO_BUFF_RD_PTR <= n55;
       end
       if ( __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ && __ILA_TX_FUNC_grant__[1] ) begin
           TXFIFO_RD_OUTPUT <= n60;
       end else if ( __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ && __ILA_TX_FUNC_grant__[2] ) begin
           TXFIFO_RD_OUTPUT <= n67;
       end
       if ( __ILA_TX_FUNC_decode_of_SET_B2B_CNTR_10G__ && __ILA_TX_FUNC_grant__[0] ) begin
           TXFIFO_RD_EN <= 1'd0;
       end
       if ( __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ && __ILA_TX_FUNC_grant__[1] ) begin
           TXFIFO_RD_EMPTY <= n71;
       end else if ( __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ && __ILA_TX_FUNC_grant__[2] ) begin
           TXFIFO_RD_EMPTY <= n75;
       end
       if ( __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ && __ILA_TX_FUNC_grant__[1] ) begin
           TX_STATE <= 5'd8;
       end else if ( __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ && __ILA_TX_FUNC_grant__[2] ) begin
           TX_STATE <= n79;
       end else if ( __ILA_TX_FUNC_decode_of_WR_PKT_LASTONE_10G__ && __ILA_TX_FUNC_grant__[3] ) begin
           TX_STATE <= 5'd1;
       end
       if ( __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ && __ILA_TX_FUNC_grant__[1] ) begin
           TX_STATE_ENCAP <= 8'd16;
       end else if ( __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ && __ILA_TX_FUNC_grant__[2] ) begin
           TX_STATE_ENCAP <= n81;
       end
       if ( __ILA_TX_FUNC_decode_of_SET_B2B_CNTR_10G__ && __ILA_TX_FUNC_grant__[0] ) begin
           TX_B2B_CNTR <= n84;
       end else if ( __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ && __ILA_TX_FUNC_grant__[1] ) begin
           TX_B2B_CNTR <= 6'd5;
       end else if ( __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ && __ILA_TX_FUNC_grant__[2] ) begin
           TX_B2B_CNTR <= n89;
       end else if ( __ILA_TX_FUNC_decode_of_WR_PKT_LASTONE_10G__ && __ILA_TX_FUNC_grant__[3] ) begin
           TX_B2B_CNTR <= n94;
       end
       if ( __ILA_TX_FUNC_decode_of_SET_B2B_CNTR_10G__ && __ILA_TX_FUNC_grant__[0] ) begin
           TX_B2B_OK <= n96;
       end else if ( __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ && __ILA_TX_FUNC_grant__[1] ) begin
           TX_B2B_OK <= 1'd0;
       end
       if ( __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ && __ILA_TX_FUNC_grant__[1] ) begin
           TX_PACKET_BYTE_CNT <= n97;
       end
       if ( __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ && __ILA_TX_FUNC_grant__[1] ) begin
           TX_WCNT <= n105;
       end else if ( __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ && __ILA_TX_FUNC_grant__[2] ) begin
           TX_WCNT <= n106;
       end
       if ( __ILA_TX_FUNC_decode_of_SET_B2B_CNTR_10G__ && __ILA_TX_FUNC_grant__[0] ) begin
           XGMII_DOUT_REG <= n108;
       end else if ( __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ && __ILA_TX_FUNC_grant__[1] ) begin
           XGMII_DOUT_REG <= n110;
       end else if ( __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ && __ILA_TX_FUNC_grant__[2] ) begin
           XGMII_DOUT_REG <= n1079;
       end
       if ( __ILA_TX_FUNC_decode_of_SET_B2B_CNTR_10G__ && __ILA_TX_FUNC_grant__[0] ) begin
           XGMII_COUT_REG <= 8'd255;
       end else if ( __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ && __ILA_TX_FUNC_grant__[1] ) begin
           XGMII_COUT_REG <= 8'd1;
       end else if ( __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ && __ILA_TX_FUNC_grant__[2] ) begin
           XGMII_COUT_REG <= n1119;
       end
       if ( __ILA_TX_FUNC_decode_of_WR_PKT_LASTONE_10G__ && __ILA_TX_FUNC_grant__[3] ) begin
           TX_PKT_SENT <= n1120;
       end
       if ( __ILA_TX_FUNC_decode_of_WR_PKT_LASTONE_10G__ && __ILA_TX_FUNC_grant__[3] ) begin
           TX_BYTE_SENT <= n1122;
       end
       if ( __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ && __ILA_TX_FUNC_grant__[1] ) begin
           CRC <= n1139;
       end else if ( __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ && __ILA_TX_FUNC_grant__[2] ) begin
           CRC <= n1002;
       end
       if ( __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ && __ILA_TX_FUNC_grant__[2] ) begin
           CRC_DAT_IN <= n1207;
       end
       if ( __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ && __ILA_TX_FUNC_grant__[1] ) begin
           CRC_IN <= n1228;
       end else if ( __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ && __ILA_TX_FUNC_grant__[2] ) begin
           CRC_IN <= n989;
       end
       if ( __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ && __ILA_TX_FUNC_grant__[1] ) begin
           TX_WCNT_INI <= n1229;
       end
       if ( __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ && __ILA_TX_FUNC_grant__[2] ) begin
           TX_BUF <= n145;
       end
       if ( __ILA_TX_FUNC_decode_of_SET_B2B_CNTR_10G__ && __ILA_TX_FUNC_grant__[0] ) begin
           TX_FUNC_INSTR <= 3'd0;
       end else if ( __ILA_TX_FUNC_decode_of_READ_BYTE_CNT_10G__ && __ILA_TX_FUNC_grant__[1] ) begin
           TX_FUNC_INSTR <= 3'd1;
       end else if ( __ILA_TX_FUNC_decode_of_WR_PKT_PAYLOAD_10G__ && __ILA_TX_FUNC_grant__[2] ) begin
           TX_FUNC_INSTR <= 3'd2;
       end else if ( __ILA_TX_FUNC_decode_of_WR_PKT_LASTONE_10G__ && __ILA_TX_FUNC_grant__[3] ) begin
           TX_FUNC_INSTR <= 3'd3;
       end
   end
end
endmodule
